`celldefine

module INV_X1_LVT (ZN, A);
output ZN;
input A;
endmodule

module OAI222_X1_LVT (ZN, A1, A2, B1, B2, C1, C2);
output ZN;
input A1, A2, B1, B2, C1, C2;
endmodule

module XNOR2_X1_LVT (ZN, A, B);
output ZN;
input A, B;
endmodule

`endcelldefine
