module openMSP430(aclk,aclk_en,dbg_freeze,dbg_i2c_sda_out,dbg_uart_txd,dco_enable,dco_wkup,dmem_addr,dmem_cen,dmem_din,dmem_wen,irq_acc,lfxt_enable,lfxt_wkup,mclk,dma_dout,dma_ready,dma_resp,per_addr,per_din,per_en,per_we,pmem_addr,pmem_cen,pmem_din,pmem_wen,puc_rst,smclk,smclk_en,cpu_en,dbg_en,dbg_i2c_addr,dbg_i2c_broadcast,dbg_i2c_scl,dbg_i2c_sda_in,dbg_uart_rxd,dco_clk,dmem_dout,irq,lfxt_clk,dma_addr,dma_din,dma_en,dma_priority,dma_we,dma_wkup,nmi,per_dout,pmem_dout,reset_n,scan_enable,scan_mode,wkup);
	 output aclk;
	 output aclk_en;
	 output dbg_freeze;
	 output dbg_i2c_sda_out;
	 output dbg_uart_txd;
	 output dco_enable;
	 output dco_wkup;
	 output [8:0]dmem_addr;
	 output dmem_cen;
	 output [15:0]dmem_din;
	 output [1:0]dmem_wen;
	 output [13:0]irq_acc;
	 output lfxt_enable;
	 output lfxt_wkup;
	 output mclk;
	 output [15:0]dma_dout;
	 output dma_ready;
	 output dma_resp;
	 output [13:0]per_addr;
	 output [15:0]per_din;
	 output per_en;
	 output [1:0]per_we;
	 output [10:0]pmem_addr;
	 output pmem_cen;
	 output [15:0]pmem_din;
	 output [1:0]pmem_wen;
	 output puc_rst;
	 output smclk;
	 output smclk_en;
	 input cpu_en;
	 input dbg_en;
	 input [6:0]dbg_i2c_addr;
	 input [6:0]dbg_i2c_broadcast;
	 input dbg_i2c_scl;
	 input dbg_i2c_sda_in;
	 input dbg_uart_rxd;
	 input dco_clk;
	 input [15:0]dmem_dout;
	 input [13:0]irq;
	 input lfxt_clk;
	 input [14:0]dma_addr;
	 input [15:0]dma_din;
	 input dma_en;
	 input dma_priority;
	 input [1:0]dma_we;
	 input dma_wkup;
	 input nmi;
	 input [15:0]per_dout;
	 input [15:0]pmem_dout;
	 input reset_n;
	 input scan_enable;
	 input scan_mode;
	 input wkup;

	 wire wdtnmies;
	 wire wdtifg;
	 wire wdt_wkup;
	 wire wdt_reset;
	 wire wdt_irq;
	 wire [15:0]per_dout_wdog;
	 wire scg1;
	 wire scg0;
	 wire pc_sw_wr;
	 wire [15:0]pc_sw;
	 wire oscoff;
	 wire [15:0]eu_mdb_out;
	 wire [1:0]eu_mb_wr;
	 wire eu_mb_en;
	 wire [15:0]eu_mab;
	 wire gie;
	 wire [15:0]dbg_reg_din;
	 wire cpuoff;
	 wire [15:0]pc_nxt;
	 wire [15:0]pc;
	 wire nmi_acc;
	 wire mclk_wkup;
	 wire mclk_enable;
	 wire mclk_dma_wkup;
	 wire mclk_dma_enable;
	 wire fe_mb_en;
	 wire [2:0]inst_type;
	 wire [15:0]inst_src;
	 wire [7:0]inst_so;
	 wire [15:0]inst_sext;
	 wire inst_mov;
	 wire [7:0]inst_jmp;
	 wire inst_irq_rst;
	 wire [15:0]inst_dext;
	 wire [15:0]inst_dest;
	 wire inst_bw;
	 wire [11:0]inst_alu;
	 wire [7:0]inst_as;
	 wire [7:0]inst_ad;
	 wire exec_done;
	 wire [3:0]e_state;
	 wire decode_noirq;
	 wire cpu_halt_st;
	 wire [15:0]per_dout_mpy;
	 wire fe_pmem_wait;
	 wire [15:0]fe_mdb_in;
	 wire [15:0]eu_mdb_in;
	 wire [15:0]dbg_mem_din;
	 wire cpu_halt_cmd;
	 wire dbg_reg_wr;
	 wire [1:0]dbg_mem_wr;
	 wire dbg_mem_en;
	 wire [15:0]dbg_mem_dout;
	 wire [15:0]dbg_mem_addr;
	 wire dbg_halt_cmd;
	 wire dbg_cpu_reset;
	 wire wdtifg_sw_set;
	 wire wdtifg_sw_clr;
	 wire wdtie;
	 wire [15:0]per_dout_sfr;
	 wire nmi_wkup;
	 wire nmi_pnd;
	 wire [31:0]cpu_id;
	 wire puc_pnd_set;
	 wire por;
	 wire [15:0]per_dout_clk;
	 wire dbg_rst;
	 wire dbg_en_s;
	 wire dbg_clk;
	 wire cpu_mclk;
	 wire cpu_en_s;
	 wire n_0_0_0;
	 wire [15:0]per_dout_or;
	 wire n_0_0_1;
	 wire n_0_0_2;
	 wire n_0_0_3;
	 wire n_0_0_4;
	 wire n_0_0_5;
	 wire n_0_0_6;
	 wire n_0_0_7;
	 wire n_0_0_8;
	 wire n_0_0_9;
	 wire n_0_0_10;
	 wire n_0_0_11;
	 wire n_0_0_12;
	 wire n_0_0_13;
	 wire n_0_0_14;
	 wire n_0_0_15;
	 wire n_14;
	 wire n_13;
	 wire n_12;
	 wire n_11;
	 wire n_10;
	 wire n_9;
	 wire n_8;
	 wire n_7;
	 wire n_6;
	 wire n_5;
	 wire n_4;
	 wire n_3;
	 wire n_2;
	 wire n_1;
	 wire n_0;
	 wire uc_0;
	 wire watchdog_0_wdt_rst_noscan;
	 wire watchdog_0_wdt_rst;
	 wire watchdog_0_wdtcnt_incr;
	 wire watchdog_0_wdtcnt_clr_sync;
	 wire watchdog_0_wdt_evt_toggle_sync;
	 wire watchdog_0_wdt_wkup_pre;
	 wire watchdog_0_n_0_0;
	 wire watchdog_0_n_0_1;
	 wire watchdog_0_n_0_2;
	 wire watchdog_0_n_0_3;
	 wire watchdog_0_n_0_4;
	 wire watchdog_0_reg_wr;
	 wire [7:0]watchdog_0_wdtctl;
	 wire watchdog_0_n_8_0;
	 wire watchdog_0_n_8_1;
	 wire watchdog_0_n_8_2;
	 wire watchdog_0_wdtpw_error;
	 wire watchdog_0_wdt_evt_toggle_sync_dly;
	 wire watchdog_0_n_9_0;
	 wire watchdog_0_wdtifg_set;
	 wire watchdog_0_n_10_0;
	 wire watchdog_0_wdtifg_clr;
	 wire watchdog_0_n_13_0;
	 wire watchdog_0_n_13_1;
	 wire watchdog_0_n_17_0;
	 wire watchdog_0_wdtcnt_clr_sync_dly;
	 wire watchdog_0_n_19_0;
	 wire watchdog_0_wdtcnt_clr;
	 wire [15:0]watchdog_0_wdtcnt;
	 wire watchdog_0_n_21_0;
	 wire watchdog_0_n_22_0;
	 wire watchdog_0_n_22_1;
	 wire [15:0]watchdog_0_wdtcnt_nxt;
	 wire watchdog_0_n_24_0;
	 wire watchdog_0_n_24_1;
	 wire watchdog_0_n_24_2;
	 wire watchdog_0_n_24_3;
	 wire watchdog_0_n_24_4;
	 wire watchdog_0_n_24_5;
	 wire watchdog_0_n_24_6;
	 wire watchdog_0_n_24_7;
	 wire watchdog_0_n_24_8;
	 wire watchdog_0_n_24_9;
	 wire watchdog_0_n_24_10;
	 wire watchdog_0_n_24_11;
	 wire watchdog_0_n_24_12;
	 wire watchdog_0_n_24_13;
	 wire watchdog_0_n_24_14;
	 wire [1:0]watchdog_0_wdtisx_ss;
	 wire [1:0]watchdog_0_wdtisx_s;
	 wire watchdog_0_n_28_0;
	 wire watchdog_0_n_28_1;
	 wire watchdog_0_n_28_2;
	 wire watchdog_0_n_28_3;
	 wire watchdog_0_n_28_4;
	 wire watchdog_0_n_28_5;
	 wire watchdog_0_n_28_6;
	 wire watchdog_0_n_28_7;
	 wire watchdog_0_n_28_8;
	 wire watchdog_0_wdtqn_reg;
	 wire watchdog_0_wdtqn_edge;
	 wire watchdog_0_wdt_evt_toggle;
	 wire watchdog_0_wdt_wkup_en;
	 wire watchdog_0_n_35_0;
	 wire watchdog_0_n_35_1;
	 wire watchdog_0_n_37_0;
	 wire watchdog_0_wdtcnt_clr_detect;
	 wire watchdog_0_wdtcnt_clr_toggle;
	 wire watchdog_0_wdtifg_clr_reg;
	 wire watchdog_0_wdtqn_edge_reg;
	 wire watchdog_0_n_1;
	 wire watchdog_0_n_0;
	 wire watchdog_0_n_2;
	 wire watchdog_0_n_3;
	 wire watchdog_0_n_4;
	 wire watchdog_0_n_30;
	 wire watchdog_0_n_29;
	 wire watchdog_0_n_35;
	 wire watchdog_0_n_34;
	 wire watchdog_0_n_17;
	 wire watchdog_0_n_31;
	 wire watchdog_0_n_33;
	 wire watchdog_0_n_27;
	 wire watchdog_0_n_10;
	 wire watchdog_0_n_16;
	 wire watchdog_0_n_15;
	 wire watchdog_0_n_14;
	 wire watchdog_0_n_13;
	 wire watchdog_0_n_12;
	 wire watchdog_0_n_11;
	 wire watchdog_0_n_26;
	 wire watchdog_0_n_25;
	 wire watchdog_0_n_24;
	 wire watchdog_0_n_23;
	 wire watchdog_0_n_22;
	 wire watchdog_0_n_21;
	 wire watchdog_0_n_20;
	 wire watchdog_0_n_19;
	 wire watchdog_0_n_18;
	 wire watchdog_0_n_28;
	 wire watchdog_0_n_7;
	 wire watchdog_0_n_5;
	 wire watchdog_0_n_6;
	 wire watchdog_0_n_8;
	 wire watchdog_0_n_9;
	 wire watchdog_0_n_32;
	 wire watchdog_0_sync_reset_por_n_0;
	 wire watchdog_0_sync_reset_por_n_1;
	 wire watchdog_0_scan_mux_wdt_rst_n_0_0;
	 wire watchdog_0_scan_mux_wdt_rst_n_0_1;
	 wire watchdog_0_sync_cell_wdtcnt_clr_n_0;
	 wire watchdog_0_sync_cell_wdtcnt_clr_n_1;
	 wire watchdog_0_sync_cell_wdtcnt_incr_n_0;
	 wire watchdog_0_sync_cell_wdtcnt_incr_n_1;
	 wire watchdog_0_sync_cell_wdt_evt_n_0;
	 wire watchdog_0_sync_cell_wdt_evt_n_1;
	 wire watchdog_0_wakeup_cell_wdog_wkup_rst;
	 wire watchdog_0_wakeup_cell_wdog_wkup_clk;
	 wire watchdog_0_wakeup_cell_wdog_n_0;
	 wire watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_0;
	 wire watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_1;
	 wire watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_0;
	 wire watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_1;
	 wire sfr_0_nmi_capture;
	 wire sfr_0_nmi_s;
	 wire sfr_0_n_0_0;
	 wire sfr_0_n_0_1;
	 wire sfr_0_n_0_2;
	 wire sfr_0_n_0_3;
	 wire sfr_0_reg_sel;
	 wire sfr_0_reg_lo_write;
	 wire sfr_0_n_2_0;
	 wire sfr_0_n_2_1;
	 wire sfr_0_n_2_2;
	 wire sfr_0_n_2_3;
	 wire sfr_0_n_2_4;
	 wire sfr_0_n_2_5;
	 wire sfr_0_n_2_6;
	 wire sfr_0_ifg1_wr;
	 wire sfr_0_nmi_capture_rst;
	 wire sfr_0_n_4_0;
	 wire sfr_0_nmie;
	 wire sfr_0_n_7_0;
	 wire sfr_0_n_8_0;
	 wire sfr_0_n_8_1;
	 wire sfr_0_nmi_dly;
	 wire sfr_0_n_10_0;
	 wire sfr_0_nmi_edge;
	 wire sfr_0_nmiifg;
	 wire sfr_0_n_13_0;
	 wire sfr_0_n_13_1;
	 wire sfr_0_n_14_0;
	 wire sfr_0_n_14_1;
	 wire sfr_0_reg_read;
	 wire sfr_0_n_27_0;
	 wire sfr_0_n_28_0;
	 wire sfr_0_nmi_pol;
	 wire sfr_0_n_1;
	 wire sfr_0_n_6;
	 wire sfr_0_n_11;
	 wire sfr_0_n_12;
	 wire sfr_0_n_13;
	 wire sfr_0_n_10;
	 wire sfr_0_n_8;
	 wire sfr_0_n_0;
	 wire sfr_0_n_5;
	 wire sfr_0_n_9;
	 wire sfr_0_n_7;
	 wire sfr_0_n_31;
	 wire sfr_0_n_14;
	 wire sfr_0_n_4;
	 wire sfr_0_n_19;
	 wire sfr_0_n_3;
	 wire sfr_0_n_18;
	 wire sfr_0_n_25;
	 wire sfr_0_n_2;
	 wire sfr_0_n_17;
	 wire sfr_0_n_24;
	 wire sfr_0_n_15;
	 wire sfr_0_n_30;
	 wire sfr_0_n_16;
	 wire sfr_0_n_27;
	 wire sfr_0_n_23;
	 wire sfr_0_n_22;
	 wire sfr_0_n_21;
	 wire sfr_0_n_26;
	 wire sfr_0_n_20;
	 wire sfr_0_n_28;
	 wire sfr_0_n_29;
	 wire sfr_0_wakeup_cell_nmi_wkup_rst;
	 wire sfr_0_wakeup_cell_nmi_wkup_clk;
	 wire sfr_0_wakeup_cell_nmi_n_0;
	 wire sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_0;
	 wire sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_1;
	 wire sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_0;
	 wire sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_1;
	 wire sfr_0_sync_cell_nmi_n_0;
	 wire sfr_0_sync_cell_nmi_n_1;
	 wire dbg_0_dbg_wr;
	 wire dbg_0_dbg_rd;
	 wire [15:0]dbg_0_dbg_din;
	 wire [5:0]dbg_0_dbg_addr;
	 wire dbg_0_n_0_0;
	 wire dbg_0_n_0_1;
	 wire dbg_0_n_0_2;
	 wire dbg_0_n_0_3;
	 wire dbg_0_mem_start;
	 wire [2:0]dbg_0_mem_ctl;
	 wire dbg_0_mem_burst_rd;
	 wire dbg_0_mem_startb;
	 wire dbg_0_n_6_0;
	 wire dbg_0_n_6_1;
	 wire dbg_0_n_8_0;
	 wire dbg_0_n_9_0;
	 wire dbg_0_n_9_1;
	 wire dbg_0_n_9_2;
	 wire dbg_0_n_9_3;
	 wire dbg_0_n_9_4;
	 wire dbg_0_n_9_5;
	 wire [1:0]dbg_0_mem_state_nxt_reg;
	 wire dbg_0_n_9_6;
	 wire [1:0]dbg_0_mem_state;
	 wire dbg_0_n_12_0;
	 wire dbg_0_mem_access;
	 wire dbg_0_n_16_0;
	 wire dbg_0_n_17_0;
	 wire dbg_0_n_17_1;
	 wire dbg_0_n_17_2;
	 wire dbg_0_n_17_3;
	 wire dbg_0_n_17_4;
	 wire dbg_0_n_17_5;
	 wire dbg_0_n_17_6;
	 wire dbg_0_n_19_0;
	 wire dbg_0_n_19_1;
	 wire dbg_0_n_19_2;
	 wire dbg_0_n_19_3;
	 wire dbg_0_n_19_4;
	 wire dbg_0_n_19_5;
	 wire dbg_0_n_19_6;
	 wire dbg_0_n_19_7;
	 wire dbg_0_n_19_8;
	 wire dbg_0_n_19_9;
	 wire dbg_0_n_19_10;
	 wire dbg_0_n_19_11;
	 wire dbg_0_n_19_12;
	 wire dbg_0_n_19_13;
	 wire dbg_0_n_19_14;
	 wire dbg_0_n_19_15;
	 wire dbg_0_n_20_0;
	 wire dbg_0_n_20_1;
	 wire dbg_0_n_20_2;
	 wire dbg_0_n_20_3;
	 wire dbg_0_n_20_4;
	 wire dbg_0_n_20_5;
	 wire dbg_0_n_20_6;
	 wire dbg_0_n_20_7;
	 wire dbg_0_n_20_8;
	 wire dbg_0_n_20_9;
	 wire dbg_0_n_20_10;
	 wire dbg_0_n_20_11;
	 wire dbg_0_n_20_12;
	 wire dbg_0_n_20_13;
	 wire dbg_0_n_20_14;
	 wire dbg_0_n_20_15;
	 wire dbg_0_n_20_16;
	 wire dbg_0_n_22_0;
	 wire dbg_0_dbg_reg_rd;
	 wire dbg_0_dbg_mem_rd;
	 wire dbg_0_dbg_mem_rd_dly;
	 wire dbg_0_dbg_rd_rdy;
	 wire dbg_0_n_32_0;
	 wire dbg_0_n_32_1;
	 wire dbg_0_n_34_0;
	 wire dbg_0_dbg_mem_acc;
	 wire dbg_0_n_35_0;
	 wire dbg_0_n_35_1;
	 wire dbg_0_n_37_0;
	 wire dbg_0_n_37_1;
	 wire dbg_0_n_37_2;
	 wire dbg_0_n_37_3;
	 wire dbg_0_n_37_4;
	 wire [15:0]dbg_0_mem_cnt;
	 wire dbg_0_n_39_0;
	 wire dbg_0_n_39_1;
	 wire dbg_0_n_39_2;
	 wire dbg_0_n_39_3;
	 wire dbg_0_n_39_4;
	 wire dbg_0_n_39_5;
	 wire dbg_0_n_39_6;
	 wire dbg_0_n_39_7;
	 wire dbg_0_n_39_8;
	 wire dbg_0_n_39_9;
	 wire dbg_0_n_39_10;
	 wire dbg_0_n_39_11;
	 wire dbg_0_n_39_12;
	 wire dbg_0_n_39_13;
	 wire dbg_0_n_39_14;
	 wire dbg_0_n_39_15;
	 wire dbg_0_n_39_16;
	 wire dbg_0_n_40_0;
	 wire dbg_0_n_40_1;
	 wire dbg_0_n_40_2;
	 wire dbg_0_n_40_3;
	 wire dbg_0_n_40_4;
	 wire dbg_0_n_40_5;
	 wire dbg_0_n_40_6;
	 wire dbg_0_n_40_7;
	 wire dbg_0_n_40_8;
	 wire dbg_0_n_40_9;
	 wire dbg_0_n_40_10;
	 wire dbg_0_n_40_11;
	 wire dbg_0_n_40_12;
	 wire dbg_0_n_40_13;
	 wire dbg_0_n_40_14;
	 wire dbg_0_n_40_15;
	 wire dbg_0_n_40_16;
	 wire dbg_0_n_42_0;
	 wire dbg_0_n_42_1;
	 wire dbg_0_n_42_2;
	 wire dbg_0_n_42_3;
	 wire dbg_0_mem_burst_start;
	 wire dbg_0_n_44_0;
	 wire dbg_0_mem_burst_end;
	 wire dbg_0_mem_burst;
	 wire dbg_0_n_46_0;
	 wire dbg_0_n_46_1;
	 wire dbg_0_n_48_0;
	 wire [5:0]dbg_0_dbg_addr_in;
	 wire dbg_0_n_48_1;
	 wire dbg_0_n_48_2;
	 wire dbg_0_n_49_0;
	 wire dbg_0_n_49_1;
	 wire dbg_0_n_49_2;
	 wire dbg_0_n_49_3;
	 wire dbg_0_n_49_4;
	 wire dbg_0_n_49_5;
	 wire dbg_0_n_49_6;
	 wire dbg_0_n_49_7;
	 wire dbg_0_n_49_8;
	 wire dbg_0_n_49_9;
	 wire dbg_0_n_49_10;
	 wire dbg_0_n_49_11;
	 wire dbg_0_n_49_12;
	 wire dbg_0_n_49_13;
	 wire dbg_0_n_49_14;
	 wire dbg_0_n_49_15;
	 wire dbg_0_n_49_16;
	 wire dbg_0_n_49_17;
	 wire dbg_0_n_49_18;
	 wire dbg_0_n_49_19;
	 wire dbg_0_n_49_20;
	 wire dbg_0_n_49_21;
	 wire dbg_0_cpu_ctl_wr;
	 wire dbg_0_mem_ctl_wr;
	 wire dbg_0_mem_data_wr;
	 wire [3:0]dbg_0_cpu_ctl;
	 wire dbg_0_n_53_0;
	 wire dbg_0_n_53_1;
	 wire dbg_0_n_54_0;
	 wire dbg_0_n_54_1;
	 wire dbg_0_n_54_2;
	 wire dbg_0_n_54_3;
	 wire dbg_0_n_54_4;
	 wire dbg_0_dbg_swbrk;
	 wire dbg_0_n_55_0;
	 wire dbg_0_n_55_1;
	 wire dbg_0_n_55_2;
	 wire dbg_0_n_55_3;
	 wire dbg_0_n_55_4;
	 wire dbg_0_n_55_5;
	 wire dbg_0_halt_flag_set;
	 wire dbg_0_n_57_0;
	 wire dbg_0_n_57_1;
	 wire dbg_0_n_57_2;
	 wire dbg_0_halt_flag_clr;
	 wire dbg_0_halt_flag;
	 wire dbg_0_n_59_0;
	 wire dbg_0_n_60_0;
	 wire dbg_0_n_60_1;
	 wire dbg_0_istep;
	 wire dbg_0_n_64_0;
	 wire dbg_0_n_64_1;
	 wire dbg_0_n_66_0;
	 wire dbg_0_n_68_0;
	 wire dbg_0_n_68_1;
	 wire dbg_0_n_68_2;
	 wire dbg_0_n_68_3;
	 wire dbg_0_n_68_4;
	 wire dbg_0_n_68_5;
	 wire dbg_0_n_68_6;
	 wire dbg_0_n_68_7;
	 wire dbg_0_n_68_8;
	 wire [15:0]dbg_0_mem_data;
	 wire dbg_0_n_70_0;
	 wire dbg_0_n_71_0;
	 wire dbg_0_n_71_1;
	 wire dbg_0_n_71_2;
	 wire dbg_0_n_71_3;
	 wire dbg_0_n_71_4;
	 wire dbg_0_n_71_5;
	 wire dbg_0_n_71_6;
	 wire dbg_0_n_71_7;
	 wire dbg_0_n_71_8;
	 wire dbg_0_n_71_9;
	 wire dbg_0_n_71_10;
	 wire dbg_0_n_71_11;
	 wire dbg_0_n_71_12;
	 wire dbg_0_n_71_13;
	 wire dbg_0_n_71_14;
	 wire dbg_0_n_71_15;
	 wire dbg_0_n_72_0;
	 wire dbg_0_n_72_1;
	 wire dbg_0_n_72_2;
	 wire dbg_0_n_74_0;
	 wire dbg_0_n_74_1;
	 wire dbg_0_n_74_2;
	 wire dbg_0_n_74_3;
	 wire dbg_0_n_74_4;
	 wire dbg_0_n_74_5;
	 wire dbg_0_n_74_6;
	 wire dbg_0_n_74_7;
	 wire dbg_0_n_74_8;
	 wire dbg_0_n_74_9;
	 wire dbg_0_n_74_10;
	 wire dbg_0_n_74_11;
	 wire dbg_0_n_74_12;
	 wire dbg_0_n_74_13;
	 wire dbg_0_n_74_14;
	 wire dbg_0_n_74_15;
	 wire dbg_0_n_74_16;
	 wire dbg_0_n_74_17;
	 wire dbg_0_n_74_18;
	 wire dbg_0_n_74_19;
	 wire [1:0]dbg_0_cpu_stat;
	 wire dbg_0_n_76_0;
	 wire dbg_0_n_76_1;
	 wire dbg_0_n_76_2;
	 wire dbg_0_n_76_3;
	 wire dbg_0_n_76_4;
	 wire dbg_0_n_76_5;
	 wire dbg_0_n_76_6;
	 wire dbg_0_n_78_0;
	 wire dbg_0_n_78_1;
	 wire dbg_0_n_78_2;
	 wire dbg_0_n_78_3;
	 wire dbg_0_n_78_4;
	 wire dbg_0_n_78_5;
	 wire dbg_0_n_78_6;
	 wire dbg_0_n_78_7;
	 wire [15:0]dbg_0_dbg_dout;
	 wire dbg_0_n_78_8;
	 wire dbg_0_n_78_9;
	 wire dbg_0_n_78_10;
	 wire dbg_0_n_78_11;
	 wire dbg_0_n_78_12;
	 wire dbg_0_n_78_13;
	 wire dbg_0_n_78_14;
	 wire dbg_0_n_78_15;
	 wire dbg_0_n_78_16;
	 wire dbg_0_n_78_17;
	 wire dbg_0_n_78_18;
	 wire dbg_0_n_78_19;
	 wire dbg_0_n_78_20;
	 wire dbg_0_n_78_21;
	 wire dbg_0_n_78_22;
	 wire dbg_0_n_78_23;
	 wire dbg_0_n_78_24;
	 wire dbg_0_n_78_25;
	 wire dbg_0_n_78_26;
	 wire dbg_0_n_78_27;
	 wire dbg_0_n_78_28;
	 wire dbg_0_n_78_29;
	 wire dbg_0_n_78_30;
	 wire dbg_0_n_78_31;
	 wire dbg_0_n_78_32;
	 wire dbg_0_n_78_33;
	 wire dbg_0_n_78_34;
	 wire dbg_0_n_78_35;
	 wire dbg_0_n_78_36;
	 wire dbg_0_n_78_37;
	 wire dbg_0_n_78_38;
	 wire dbg_0_n_78_39;
	 wire dbg_0_n_78_40;
	 wire dbg_0_n_78_41;
	 wire dbg_0_n_78_42;
	 wire dbg_0_n_78_43;
	 wire dbg_0_n_78_44;
	 wire dbg_0_n_78_45;
	 wire dbg_0_n_78_46;
	 wire dbg_0_n_78_47;
	 wire dbg_0_n_78_48;
	 wire dbg_0_n_78_49;
	 wire dbg_0_n_78_50;
	 wire dbg_0_n_78_51;
	 wire dbg_0_n_78_52;
	 wire dbg_0_n_78_53;
	 wire dbg_0_n_78_54;
	 wire dbg_0_n_78_55;
	 wire dbg_0_n_78_56;
	 wire dbg_0_n_78_57;
	 wire dbg_0_n_78_58;
	 wire dbg_0_n_78_59;
	 wire dbg_0_n_78_60;
	 wire dbg_0_n_78_61;
	 wire dbg_0_n_78_62;
	 wire dbg_0_n_78_63;
	 wire dbg_0_n_78_64;
	 wire dbg_0_n_78_65;
	 wire dbg_0_n_78_66;
	 wire dbg_0_n_78_67;
	 wire dbg_0_n_78_68;
	 wire dbg_0_n_78_69;
	 wire dbg_0_n_78_70;
	 wire dbg_0_n_78_71;
	 wire dbg_0_n_78_72;
	 wire dbg_0_n_78_73;
	 wire dbg_0_n_78_74;
	 wire dbg_0_n_78_75;
	 wire dbg_0_n_78_76;
	 wire dbg_0_n_78_77;
	 wire dbg_0_n_78_78;
	 wire dbg_0_n_78_79;
	 wire dbg_0_n_78_80;
	 wire dbg_0_n_78_81;
	 wire dbg_0_n_78_82;
	 wire dbg_0_n_78_83;
	 wire dbg_0_n_78_84;
	 wire dbg_0_n_78_85;
	 wire dbg_0_n_78_86;
	 wire dbg_0_n_78_87;
	 wire dbg_0_n_78_88;
	 wire dbg_0_n_78_89;
	 wire dbg_0_n_78_90;
	 wire dbg_0_n_78_91;
	 wire dbg_0_n_78_92;
	 wire dbg_0_n_78_93;
	 wire dbg_0_n_78_94;
	 wire dbg_0_n_78_95;
	 wire dbg_0_n_78_96;
	 wire dbg_0_n_78_97;
	 wire dbg_0_n_78_98;
	 wire dbg_0_n_78_99;
	 wire dbg_0_n_78_100;
	 wire dbg_0_n_78_101;
	 wire dbg_0_n_78_102;
	 wire dbg_0_n_78_103;
	 wire dbg_0_n_78_104;
	 wire dbg_0_n_78_105;
	 wire dbg_0_n_78_106;
	 wire dbg_0_n_78_107;
	 wire dbg_0_n_78_108;
	 wire dbg_0_n_78_109;
	 wire dbg_0_n_78_110;
	 wire dbg_0_n_78_111;
	 wire dbg_0_n_78_112;
	 wire dbg_0_n_78_113;
	 wire dbg_0_n_78_114;
	 wire dbg_0_n_78_115;
	 wire dbg_0_mem_burst_wr;
	 wire dbg_0_n_95;
	 wire dbg_0_n_1;
	 wire dbg_0_n_104;
	 wire dbg_0_n_98;
	 wire dbg_0_n_102;
	 wire dbg_0_n_55;
	 wire dbg_0_n_57;
	 wire dbg_0_n_73;
	 wire dbg_0_n_58;
	 wire dbg_0_n_74;
	 wire dbg_0_n_59;
	 wire dbg_0_n_75;
	 wire dbg_0_n_60;
	 wire dbg_0_n_76;
	 wire dbg_0_n_61;
	 wire dbg_0_n_77;
	 wire dbg_0_n_62;
	 wire dbg_0_n_78;
	 wire dbg_0_n_63;
	 wire dbg_0_n_79;
	 wire dbg_0_n_64;
	 wire dbg_0_n_80;
	 wire dbg_0_n_65;
	 wire dbg_0_n_81;
	 wire dbg_0_n_66;
	 wire dbg_0_n_82;
	 wire dbg_0_n_67;
	 wire dbg_0_n_83;
	 wire dbg_0_n_68;
	 wire dbg_0_n_84;
	 wire dbg_0_n_69;
	 wire dbg_0_n_85;
	 wire dbg_0_n_70;
	 wire dbg_0_n_86;
	 wire dbg_0_n_71;
	 wire dbg_0_n_87;
	 wire dbg_0_n_2;
	 wire dbg_0_n_3;
	 wire dbg_0_n_4;
	 wire dbg_0_n_0;
	 wire dbg_0_n_5;
	 wire dbg_0_n_6;
	 wire dbg_0_n_7;
	 wire dbg_0_n_47;
	 wire dbg_0_n_48;
	 wire dbg_0_n_96;
	 wire dbg_0_n_101;
	 wire dbg_0_n_10;
	 wire dbg_0_n_53;
	 wire dbg_0_n_11;
	 wire dbg_0_n_13;
	 wire dbg_0_n_29;
	 wire dbg_0_n_46;
	 wire dbg_0_n_45;
	 wire dbg_0_n_49;
	 wire dbg_0_n_51;
	 wire dbg_0_n_9;
	 wire dbg_0_n_50;
	 wire dbg_0_n_52;
	 wire dbg_0_n_54;
	 wire dbg_0_n_56;
	 wire dbg_0_n_72;
	 wire dbg_0_n_88;
	 wire dbg_0_n_90;
	 wire dbg_0_n_89;
	 wire dbg_0_n_27;
	 wire dbg_0_n_43;
	 wire dbg_0_n_26;
	 wire dbg_0_n_42;
	 wire dbg_0_n_25;
	 wire dbg_0_n_41;
	 wire dbg_0_n_24;
	 wire dbg_0_n_40;
	 wire dbg_0_n_23;
	 wire dbg_0_n_39;
	 wire dbg_0_n_22;
	 wire dbg_0_n_38;
	 wire dbg_0_n_21;
	 wire dbg_0_n_37;
	 wire dbg_0_n_20;
	 wire dbg_0_n_36;
	 wire dbg_0_n_19;
	 wire dbg_0_n_35;
	 wire dbg_0_n_18;
	 wire dbg_0_n_34;
	 wire dbg_0_n_17;
	 wire dbg_0_n_33;
	 wire dbg_0_n_16;
	 wire dbg_0_n_32;
	 wire dbg_0_n_15;
	 wire dbg_0_n_31;
	 wire dbg_0_n_12;
	 wire dbg_0_n_14;
	 wire dbg_0_n_30;
	 wire dbg_0_n_28;
	 wire dbg_0_n_44;
	 wire dbg_0_n_97;
	 wire dbg_0_n_136;
	 wire dbg_0_n_135;
	 wire dbg_0_n_115;
	 wire dbg_0_n_133;
	 wire dbg_0_n_152;
	 wire dbg_0_n_153;
	 wire dbg_0_n_134;
	 wire dbg_0_n_92;
	 wire dbg_0_n_91;
	 wire dbg_0_n_99;
	 wire dbg_0_n_132;
	 wire dbg_0_n_151;
	 wire dbg_0_n_131;
	 wire dbg_0_n_150;
	 wire dbg_0_n_130;
	 wire dbg_0_n_149;
	 wire dbg_0_n_129;
	 wire dbg_0_n_148;
	 wire dbg_0_n_128;
	 wire dbg_0_n_147;
	 wire dbg_0_n_127;
	 wire dbg_0_n_146;
	 wire dbg_0_n_126;
	 wire dbg_0_n_145;
	 wire dbg_0_n_116;
	 wire dbg_0_n_117;
	 wire dbg_0_n_125;
	 wire dbg_0_n_144;
	 wire dbg_0_n_124;
	 wire dbg_0_n_143;
	 wire dbg_0_n_93;
	 wire dbg_0_n_123;
	 wire dbg_0_n_142;
	 wire dbg_0_n_105;
	 wire dbg_0_n_122;
	 wire dbg_0_n_141;
	 wire dbg_0_n_106;
	 wire dbg_0_n_121;
	 wire dbg_0_n_140;
	 wire dbg_0_n_94;
	 wire dbg_0_n_107;
	 wire dbg_0_n_100;
	 wire dbg_0_n_155;
	 wire dbg_0_n_120;
	 wire dbg_0_n_139;
	 wire dbg_0_n_154;
	 wire dbg_0_n_119;
	 wire dbg_0_n_138;
	 wire dbg_0_n_118;
	 wire dbg_0_n_137;
	 wire dbg_0_n_103;
	 wire dbg_0_n_8;
	 wire dbg_0_n_108;
	 wire dbg_0_n_110;
	 wire dbg_0_n_111;
	 wire dbg_0_n_109;
	 wire dbg_0_n_113;
	 wire dbg_0_n_114;
	 wire dbg_0_n_112;
	 wire dbg_0_dbg_uart_0_uart_rxd_n;
	 wire dbg_0_dbg_uart_0_uart_rxd;
	 wire [1:0]dbg_0_dbg_uart_0_rxd_buf;
	 wire dbg_0_dbg_uart_0_n_2_0;
	 wire dbg_0_dbg_uart_0_n_2_1;
	 wire dbg_0_dbg_uart_0_n_2_2;
	 wire dbg_0_dbg_uart_0_rxd_maj_nxt;
	 wire [19:0]dbg_0_dbg_uart_0_xfer_buf;
	 wire dbg_0_dbg_uart_0_n_4_0;
	 wire dbg_0_dbg_uart_0_n_4_1;
	 wire dbg_0_dbg_uart_0_n_4_2;
	 wire dbg_0_dbg_uart_0_n_4_3;
	 wire dbg_0_dbg_uart_0_n_4_4;
	 wire dbg_0_dbg_uart_0_n_4_5;
	 wire dbg_0_dbg_uart_0_n_4_6;
	 wire dbg_0_dbg_uart_0_n_4_7;
	 wire dbg_0_dbg_uart_0_n_4_8;
	 wire dbg_0_dbg_uart_0_n_4_9;
	 wire dbg_0_dbg_uart_0_n_4_10;
	 wire dbg_0_dbg_uart_0_n_4_11;
	 wire dbg_0_dbg_uart_0_n_4_12;
	 wire dbg_0_dbg_uart_0_n_4_13;
	 wire dbg_0_dbg_uart_0_n_4_14;
	 wire dbg_0_dbg_uart_0_n_4_15;
	 wire dbg_0_dbg_uart_0_n_4_16;
	 wire dbg_0_dbg_uart_0_n_4_17;
	 wire dbg_0_dbg_uart_0_n_4_18;
	 wire dbg_0_dbg_uart_0_n_5_0;
	 wire dbg_0_dbg_uart_0_n_5_1;
	 wire dbg_0_dbg_uart_0_rxd_maj;
	 wire dbg_0_dbg_uart_0_n_7_0;
	 wire dbg_0_dbg_uart_0_n_8_0;
	 wire dbg_0_dbg_uart_0_n_8_1;
	 wire dbg_0_dbg_uart_0_n_8_2;
	 wire dbg_0_dbg_uart_0_n_8_3;
	 wire dbg_0_dbg_uart_0_n_8_4;
	 wire dbg_0_dbg_uart_0_n_8_5;
	 wire dbg_0_dbg_uart_0_n_8_6;
	 wire dbg_0_dbg_uart_0_n_8_7;
	 wire dbg_0_dbg_uart_0_n_8_8;
	 wire dbg_0_dbg_uart_0_n_8_9;
	 wire dbg_0_dbg_uart_0_n_8_10;
	 wire dbg_0_dbg_uart_0_n_8_11;
	 wire dbg_0_dbg_uart_0_n_8_12;
	 wire dbg_0_dbg_uart_0_n_8_13;
	 wire dbg_0_dbg_uart_0_n_8_14;
	 wire dbg_0_dbg_uart_0_n_8_15;
	 wire dbg_0_dbg_uart_0_n_8_16;
	 wire dbg_0_dbg_uart_0_n_8_17;
	 wire dbg_0_dbg_uart_0_n_8_18;
	 wire dbg_0_dbg_uart_0_n_8_19;
	 wire dbg_0_dbg_uart_0_n_8_20;
	 wire dbg_0_dbg_uart_0_n_8_21;
	 wire dbg_0_dbg_uart_0_n_8_22;
	 wire dbg_0_dbg_uart_0_n_8_23;
	 wire dbg_0_dbg_uart_0_n_8_24;
	 wire [2:0]dbg_0_dbg_uart_0_uart_state_nxt_reg;
	 wire dbg_0_dbg_uart_0_n_8_25;
	 wire dbg_0_dbg_uart_0_n_8_26;
	 wire dbg_0_dbg_uart_0_n_8_27;
	 wire dbg_0_dbg_uart_0_n_8_28;
	 wire dbg_0_dbg_uart_0_n_8_29;
	 wire [2:0]dbg_0_dbg_uart_0_uart_state;
	 wire dbg_0_dbg_uart_0_n_11_0;
	 wire dbg_0_dbg_uart_0_n_11_1;
	 wire dbg_0_dbg_uart_0_n_13_0;
	 wire dbg_0_dbg_uart_0_n_13_1;
	 wire dbg_0_dbg_uart_0_n_13_2;
	 wire dbg_0_dbg_uart_0_n_14_0;
	 wire dbg_0_dbg_uart_0_n_15_0;
	 wire dbg_0_dbg_uart_0_rxd_fe;
	 wire dbg_0_dbg_uart_0_sync_busy;
	 wire [15:0]dbg_0_dbg_uart_0_bit_cnt_max;
	 wire dbg_0_dbg_uart_0_n_21_0;
	 wire dbg_0_dbg_uart_0_n_21_1;
	 wire dbg_0_dbg_uart_0_n_21_2;
	 wire dbg_0_dbg_uart_0_n_21_3;
	 wire dbg_0_dbg_uart_0_n_21_4;
	 wire dbg_0_dbg_uart_0_n_21_5;
	 wire dbg_0_dbg_uart_0_n_21_6;
	 wire dbg_0_dbg_uart_0_n_21_7;
	 wire dbg_0_dbg_uart_0_n_21_8;
	 wire dbg_0_dbg_uart_0_n_21_9;
	 wire dbg_0_dbg_uart_0_n_21_10;
	 wire dbg_0_dbg_uart_0_n_21_11;
	 wire dbg_0_dbg_uart_0_n_21_12;
	 wire dbg_0_dbg_uart_0_n_21_13;
	 wire dbg_0_dbg_uart_0_n_21_14;
	 wire dbg_0_dbg_uart_0_n_21_15;
	 wire dbg_0_dbg_uart_0_n_21_16;
	 wire dbg_0_dbg_uart_0_n_21_17;
	 wire dbg_0_dbg_uart_0_n_22_0;
	 wire dbg_0_dbg_uart_0_n_22_1;
	 wire dbg_0_dbg_uart_0_n_24_0;
	 wire dbg_0_dbg_uart_0_txd_start;
	 wire dbg_0_dbg_uart_0_rx_active;
	 wire [15:0]dbg_0_dbg_uart_0_xfer_cnt;
	 wire dbg_0_dbg_uart_0_n_27_0;
	 wire dbg_0_dbg_uart_0_n_27_1;
	 wire dbg_0_dbg_uart_0_n_27_2;
	 wire dbg_0_dbg_uart_0_n_27_3;
	 wire dbg_0_dbg_uart_0_n_27_4;
	 wire dbg_0_dbg_uart_0_n_27_5;
	 wire dbg_0_dbg_uart_0_n_27_6;
	 wire dbg_0_dbg_uart_0_n_27_7;
	 wire dbg_0_dbg_uart_0_n_27_8;
	 wire dbg_0_dbg_uart_0_n_27_9;
	 wire dbg_0_dbg_uart_0_n_27_10;
	 wire dbg_0_dbg_uart_0_n_27_11;
	 wire dbg_0_dbg_uart_0_n_27_12;
	 wire dbg_0_dbg_uart_0_n_27_13;
	 wire dbg_0_dbg_uart_0_n_29_0;
	 wire dbg_0_dbg_uart_0_n_30_0;
	 wire dbg_0_dbg_uart_0_n_31_0;
	 wire dbg_0_dbg_uart_0_n_31_1;
	 wire dbg_0_dbg_uart_0_n_31_2;
	 wire dbg_0_dbg_uart_0_n_31_3;
	 wire dbg_0_dbg_uart_0_n_31_4;
	 wire dbg_0_dbg_uart_0_n_31_5;
	 wire dbg_0_dbg_uart_0_n_31_6;
	 wire dbg_0_dbg_uart_0_n_31_7;
	 wire dbg_0_dbg_uart_0_n_31_8;
	 wire dbg_0_dbg_uart_0_n_31_9;
	 wire dbg_0_dbg_uart_0_n_31_10;
	 wire dbg_0_dbg_uart_0_n_31_11;
	 wire dbg_0_dbg_uart_0_n_31_12;
	 wire dbg_0_dbg_uart_0_n_31_13;
	 wire dbg_0_dbg_uart_0_n_31_14;
	 wire dbg_0_dbg_uart_0_n_31_15;
	 wire dbg_0_dbg_uart_0_n_31_16;
	 wire dbg_0_dbg_uart_0_n_31_17;
	 wire dbg_0_dbg_uart_0_n_31_18;
	 wire dbg_0_dbg_uart_0_n_31_19;
	 wire dbg_0_dbg_uart_0_n_31_20;
	 wire dbg_0_dbg_uart_0_n_31_21;
	 wire dbg_0_dbg_uart_0_n_31_22;
	 wire dbg_0_dbg_uart_0_n_31_23;
	 wire dbg_0_dbg_uart_0_n_31_24;
	 wire dbg_0_dbg_uart_0_n_31_25;
	 wire dbg_0_dbg_uart_0_n_31_26;
	 wire dbg_0_dbg_uart_0_n_31_27;
	 wire dbg_0_dbg_uart_0_n_31_28;
	 wire dbg_0_dbg_uart_0_n_31_29;
	 wire dbg_0_dbg_uart_0_n_31_30;
	 wire dbg_0_dbg_uart_0_n_31_31;
	 wire dbg_0_dbg_uart_0_n_31_32;
	 wire dbg_0_dbg_uart_0_n_32_0;
	 wire dbg_0_dbg_uart_0_n_32_1;
	 wire dbg_0_dbg_uart_0_n_32_2;
	 wire dbg_0_dbg_uart_0_n_32_3;
	 wire dbg_0_dbg_uart_0_n_33_0;
	 wire dbg_0_dbg_uart_0_n_33_1;
	 wire dbg_0_dbg_uart_0_n_33_2;
	 wire dbg_0_dbg_uart_0_n_35_0;
	 wire dbg_0_dbg_uart_0_n_35_1;
	 wire dbg_0_dbg_uart_0_n_35_2;
	 wire dbg_0_dbg_uart_0_n_35_3;
	 wire dbg_0_dbg_uart_0_n_35_4;
	 wire dbg_0_dbg_uart_0_n_35_5;
	 wire dbg_0_dbg_uart_0_xfer_bit_inc;
	 wire [3:0]dbg_0_dbg_uart_0_xfer_bit;
	 wire dbg_0_dbg_uart_0_n_39_0;
	 wire dbg_0_dbg_uart_0_n_39_1;
	 wire dbg_0_dbg_uart_0_n_39_2;
	 wire dbg_0_dbg_uart_0_n_40_0;
	 wire dbg_0_dbg_uart_0_n_41_0;
	 wire dbg_0_dbg_uart_0_n_41_1;
	 wire dbg_0_dbg_uart_0_n_42_0;
	 wire dbg_0_dbg_uart_0_n_42_1;
	 wire dbg_0_dbg_uart_0_n_42_2;
	 wire dbg_0_dbg_uart_0_n_44_0;
	 wire dbg_0_dbg_uart_0_n_44_1;
	 wire dbg_0_dbg_uart_0_n_44_2;
	 wire dbg_0_dbg_uart_0_n_44_3;
	 wire dbg_0_dbg_uart_0_xfer_done;
	 wire dbg_0_dbg_uart_0_cmd_valid;
	 wire dbg_0_dbg_uart_0_dbg_bw;
	 wire dbg_0_dbg_uart_0_n_49_0;
	 wire dbg_0_dbg_uart_0_n_49_1;
	 wire dbg_0_dbg_uart_0_n_49_2;
	 wire dbg_0_dbg_uart_0_n_49_3;
	 wire dbg_0_dbg_uart_0_n_49_4;
	 wire dbg_0_dbg_uart_0_n_49_5;
	 wire dbg_0_dbg_uart_0_n_49_6;
	 wire dbg_0_dbg_uart_0_n_49_7;
	 wire dbg_0_dbg_uart_0_n_49_8;
	 wire dbg_0_dbg_uart_0_n_49_9;
	 wire dbg_0_dbg_uart_0_n_49_10;
	 wire dbg_0_dbg_uart_0_n_50_0;
	 wire dbg_0_dbg_uart_0_n_50_1;
	 wire dbg_0_dbg_uart_0_n_52_0;
	 wire dbg_0_dbg_uart_0_n_52_1;
	 wire dbg_0_dbg_uart_0_n_54_0;
	 wire dbg_0_dbg_uart_0_n_136;
	 wire dbg_0_dbg_uart_0_n_130;
	 wire dbg_0_dbg_uart_0_n_19;
	 wire dbg_0_dbg_uart_0_n_76;
	 wire dbg_0_dbg_uart_0_n_53;
	 wire dbg_0_dbg_uart_0_n_58;
	 wire dbg_0_dbg_uart_0_n_54;
	 wire dbg_0_dbg_uart_0_n_56;
	 wire dbg_0_dbg_uart_0_n_57;
	 wire dbg_0_dbg_uart_0_n_55;
	 wire dbg_0_dbg_uart_0_n_52;
	 wire dbg_0_dbg_uart_0_n_59;
	 wire dbg_0_dbg_uart_0_n_51;
	 wire dbg_0_dbg_uart_0_n_22;
	 wire dbg_0_dbg_uart_0_n_119;
	 wire dbg_0_dbg_uart_0_n_123;
	 wire dbg_0_dbg_uart_0_n_124;
	 wire dbg_0_dbg_uart_0_n_128;
	 wire dbg_0_dbg_uart_0_n_118;
	 wire dbg_0_dbg_uart_0_n_120;
	 wire dbg_0_dbg_uart_0_n_125;
	 wire dbg_0_dbg_uart_0_n_121;
	 wire dbg_0_dbg_uart_0_n_122;
	 wire dbg_0_dbg_uart_0_n_127;
	 wire dbg_0_dbg_uart_0_n_116;
	 wire dbg_0_dbg_uart_0_n_117;
	 wire dbg_0_dbg_uart_0_n_28;
	 wire dbg_0_dbg_uart_0_n_126;
	 wire dbg_0_dbg_uart_0_n_25;
	 wire dbg_0_dbg_uart_0_n_27;
	 wire dbg_0_dbg_uart_0_n_26;
	 wire dbg_0_dbg_uart_0_n_29;
	 wire dbg_0_dbg_uart_0_n_31;
	 wire dbg_0_dbg_uart_0_n_24;
	 wire dbg_0_dbg_uart_0_n_23;
	 wire dbg_0_dbg_uart_0_n_33;
	 wire dbg_0_dbg_uart_0_n_34;
	 wire dbg_0_dbg_uart_0_n_32;
	 wire dbg_0_dbg_uart_0_n_50;
	 wire dbg_0_dbg_uart_0_n_60;
	 wire dbg_0_dbg_uart_0_n_61;
	 wire dbg_0_dbg_uart_0_n_49;
	 wire dbg_0_dbg_uart_0_n_95;
	 wire dbg_0_dbg_uart_0_n_94;
	 wire dbg_0_dbg_uart_0_n_97;
	 wire dbg_0_dbg_uart_0_n_78;
	 wire dbg_0_dbg_uart_0_n_96;
	 wire dbg_0_dbg_uart_0_n_98;
	 wire dbg_0_dbg_uart_0_n_79;
	 wire dbg_0_dbg_uart_0_n_62;
	 wire dbg_0_dbg_uart_0_n_48;
	 wire dbg_0_dbg_uart_0_n_99;
	 wire dbg_0_dbg_uart_0_n_77;
	 wire dbg_0_dbg_uart_0_n_80;
	 wire dbg_0_dbg_uart_0_n_63;
	 wire dbg_0_dbg_uart_0_n_47;
	 wire dbg_0_dbg_uart_0_n_100;
	 wire dbg_0_dbg_uart_0_n_81;
	 wire dbg_0_dbg_uart_0_n_64;
	 wire dbg_0_dbg_uart_0_n_46;
	 wire dbg_0_dbg_uart_0_n_101;
	 wire dbg_0_dbg_uart_0_n_82;
	 wire dbg_0_dbg_uart_0_n_65;
	 wire dbg_0_dbg_uart_0_n_45;
	 wire dbg_0_dbg_uart_0_n_102;
	 wire dbg_0_dbg_uart_0_n_83;
	 wire dbg_0_dbg_uart_0_n_66;
	 wire dbg_0_dbg_uart_0_n_44;
	 wire dbg_0_dbg_uart_0_n_103;
	 wire dbg_0_dbg_uart_0_n_84;
	 wire dbg_0_dbg_uart_0_n_67;
	 wire dbg_0_dbg_uart_0_n_43;
	 wire dbg_0_dbg_uart_0_n_104;
	 wire dbg_0_dbg_uart_0_n_85;
	 wire dbg_0_dbg_uart_0_n_68;
	 wire dbg_0_dbg_uart_0_n_42;
	 wire dbg_0_dbg_uart_0_n_105;
	 wire dbg_0_dbg_uart_0_n_86;
	 wire dbg_0_dbg_uart_0_n_69;
	 wire dbg_0_dbg_uart_0_n_41;
	 wire dbg_0_dbg_uart_0_n_106;
	 wire dbg_0_dbg_uart_0_n_87;
	 wire dbg_0_dbg_uart_0_n_70;
	 wire dbg_0_dbg_uart_0_n_40;
	 wire dbg_0_dbg_uart_0_n_107;
	 wire dbg_0_dbg_uart_0_n_88;
	 wire dbg_0_dbg_uart_0_n_71;
	 wire dbg_0_dbg_uart_0_n_39;
	 wire dbg_0_dbg_uart_0_n_108;
	 wire dbg_0_dbg_uart_0_n_89;
	 wire dbg_0_dbg_uart_0_n_72;
	 wire dbg_0_dbg_uart_0_n_38;
	 wire dbg_0_dbg_uart_0_n_109;
	 wire dbg_0_dbg_uart_0_n_90;
	 wire dbg_0_dbg_uart_0_n_73;
	 wire dbg_0_dbg_uart_0_n_37;
	 wire dbg_0_dbg_uart_0_n_110;
	 wire dbg_0_dbg_uart_0_n_91;
	 wire dbg_0_dbg_uart_0_n_74;
	 wire dbg_0_dbg_uart_0_n_36;
	 wire dbg_0_dbg_uart_0_n_111;
	 wire dbg_0_dbg_uart_0_n_92;
	 wire dbg_0_dbg_uart_0_n_75;
	 wire dbg_0_dbg_uart_0_n_35;
	 wire dbg_0_dbg_uart_0_n_112;
	 wire dbg_0_dbg_uart_0_n_93;
	 wire dbg_0_dbg_uart_0_n_113;
	 wire dbg_0_dbg_uart_0_n_114;
	 wire dbg_0_dbg_uart_0_n_115;
	 wire dbg_0_dbg_uart_0_n_21;
	 wire dbg_0_dbg_uart_0_n_0;
	 wire dbg_0_dbg_uart_0_n_18;
	 wire dbg_0_dbg_uart_0_n_17;
	 wire dbg_0_dbg_uart_0_n_129;
	 wire dbg_0_dbg_uart_0_n_16;
	 wire dbg_0_dbg_uart_0_n_15;
	 wire dbg_0_dbg_uart_0_n_14;
	 wire dbg_0_dbg_uart_0_n_13;
	 wire dbg_0_dbg_uart_0_n_12;
	 wire dbg_0_dbg_uart_0_n_131;
	 wire dbg_0_dbg_uart_0_n_11;
	 wire dbg_0_dbg_uart_0_n_10;
	 wire dbg_0_dbg_uart_0_n_20;
	 wire dbg_0_dbg_uart_0_n_9;
	 wire dbg_0_dbg_uart_0_n_8;
	 wire dbg_0_dbg_uart_0_n_7;
	 wire dbg_0_dbg_uart_0_n_6;
	 wire dbg_0_dbg_uart_0_n_5;
	 wire dbg_0_dbg_uart_0_n_4;
	 wire dbg_0_dbg_uart_0_n_132;
	 wire dbg_0_dbg_uart_0_n_30;
	 wire dbg_0_dbg_uart_0_n_133;
	 wire dbg_0_dbg_uart_0_n_3;
	 wire dbg_0_dbg_uart_0_n_2;
	 wire dbg_0_dbg_uart_0_n_1;
	 wire dbg_0_dbg_uart_0_n_135;
	 wire dbg_0_dbg_uart_0_n_134;
	 wire dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_0;
	 wire dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_1;
	 wire multiplier_0_n_0_0;
	 wire multiplier_0_n_0_1;
	 wire multiplier_0_n_0_2;
	 wire multiplier_0_n_0_3;
	 wire multiplier_0_reg_sel;
	 wire multiplier_0_reg_read;
	 wire multiplier_0_n_3_0;
	 wire multiplier_0_n_3_1;
	 wire multiplier_0_n_3_2;
	 wire multiplier_0_reg_rd1;
	 wire multiplier_0_reg_rd15;
	 wire multiplier_0_reg_write;
	 wire multiplier_0_op2_wr;
	 wire multiplier_0_reslo_wr;
	 wire multiplier_0_reshi_wr;
	 wire [15:0]multiplier_0_per_din_msk;
	 wire [15:0]multiplier_0_op2_reg;
	 wire [1:0]multiplier_0_cycle;
	 wire multiplier_0_result_wr;
	 wire multiplier_0_op1_wr;
	 wire multiplier_0_sign_sel;
	 wire [8:0]multiplier_0_op2_hi_xp;
	 wire multiplier_0_n_29_0;
	 wire multiplier_0_n_29_1;
	 wire [8:0]multiplier_0_op2_xp;
	 wire multiplier_0_n_29_2;
	 wire multiplier_0_n_29_3;
	 wire multiplier_0_n_29_4;
	 wire multiplier_0_n_29_5;
	 wire multiplier_0_n_29_6;
	 wire multiplier_0_n_29_7;
	 wire multiplier_0_n_29_8;
	 wire [15:0]multiplier_0_op1;
	 wire [16:0]multiplier_0_op1_xp;
	 wire multiplier_0_n_32_0;
	 wire multiplier_0_n_32_1;
	 wire multiplier_0_n_32_2;
	 wire multiplier_0_n_32_3;
	 wire multiplier_0_n_32_4;
	 wire multiplier_0_n_32_5;
	 wire multiplier_0_n_32_6;
	 wire multiplier_0_n_32_7;
	 wire multiplier_0_n_32_8;
	 wire multiplier_0_n_32_9;
	 wire multiplier_0_n_32_10;
	 wire multiplier_0_n_32_11;
	 wire multiplier_0_n_32_12;
	 wire multiplier_0_n_32_13;
	 wire multiplier_0_n_32_14;
	 wire multiplier_0_n_32_15;
	 wire multiplier_0_n_32_16;
	 wire multiplier_0_n_32_17;
	 wire multiplier_0_n_32_18;
	 wire multiplier_0_n_32_19;
	 wire multiplier_0_n_32_20;
	 wire multiplier_0_n_32_21;
	 wire multiplier_0_n_32_22;
	 wire multiplier_0_n_32_23;
	 wire multiplier_0_n_32_24;
	 wire multiplier_0_n_32_25;
	 wire multiplier_0_n_32_26;
	 wire multiplier_0_n_32_27;
	 wire multiplier_0_n_32_28;
	 wire multiplier_0_n_32_29;
	 wire multiplier_0_n_32_30;
	 wire multiplier_0_n_32_31;
	 wire multiplier_0_n_32_32;
	 wire multiplier_0_n_32_33;
	 wire multiplier_0_n_32_34;
	 wire multiplier_0_n_32_35;
	 wire multiplier_0_n_32_36;
	 wire multiplier_0_n_32_37;
	 wire multiplier_0_n_32_38;
	 wire multiplier_0_n_32_39;
	 wire multiplier_0_n_32_40;
	 wire multiplier_0_n_32_41;
	 wire multiplier_0_n_32_42;
	 wire multiplier_0_n_32_43;
	 wire multiplier_0_n_32_44;
	 wire multiplier_0_n_32_45;
	 wire multiplier_0_n_32_46;
	 wire multiplier_0_n_32_47;
	 wire multiplier_0_n_32_48;
	 wire multiplier_0_n_32_49;
	 wire multiplier_0_n_32_50;
	 wire multiplier_0_n_32_51;
	 wire multiplier_0_n_32_52;
	 wire multiplier_0_n_32_53;
	 wire multiplier_0_n_32_54;
	 wire multiplier_0_n_32_55;
	 wire multiplier_0_n_32_56;
	 wire multiplier_0_n_32_57;
	 wire multiplier_0_n_32_58;
	 wire multiplier_0_n_32_59;
	 wire multiplier_0_n_32_60;
	 wire multiplier_0_n_32_61;
	 wire multiplier_0_n_32_62;
	 wire multiplier_0_n_32_63;
	 wire multiplier_0_n_32_64;
	 wire multiplier_0_n_32_65;
	 wire multiplier_0_n_32_66;
	 wire multiplier_0_n_32_67;
	 wire multiplier_0_n_32_68;
	 wire multiplier_0_n_32_69;
	 wire multiplier_0_n_32_70;
	 wire multiplier_0_n_32_71;
	 wire multiplier_0_n_32_72;
	 wire multiplier_0_n_32_73;
	 wire multiplier_0_n_32_74;
	 wire multiplier_0_n_32_75;
	 wire multiplier_0_n_32_76;
	 wire multiplier_0_n_32_77;
	 wire multiplier_0_n_32_78;
	 wire multiplier_0_n_32_79;
	 wire multiplier_0_n_32_80;
	 wire multiplier_0_n_32_81;
	 wire multiplier_0_n_32_82;
	 wire multiplier_0_n_32_83;
	 wire multiplier_0_n_32_84;
	 wire multiplier_0_n_32_85;
	 wire multiplier_0_n_32_86;
	 wire multiplier_0_n_32_87;
	 wire multiplier_0_n_32_88;
	 wire multiplier_0_n_32_89;
	 wire multiplier_0_n_32_90;
	 wire multiplier_0_n_32_91;
	 wire multiplier_0_n_32_92;
	 wire multiplier_0_n_32_93;
	 wire multiplier_0_n_32_94;
	 wire multiplier_0_n_32_95;
	 wire multiplier_0_n_32_96;
	 wire multiplier_0_n_32_97;
	 wire multiplier_0_n_32_98;
	 wire multiplier_0_n_32_99;
	 wire multiplier_0_n_32_100;
	 wire multiplier_0_n_32_101;
	 wire multiplier_0_n_32_102;
	 wire multiplier_0_n_32_103;
	 wire multiplier_0_n_32_104;
	 wire multiplier_0_n_32_105;
	 wire multiplier_0_n_32_106;
	 wire multiplier_0_n_32_107;
	 wire multiplier_0_n_32_108;
	 wire multiplier_0_n_32_109;
	 wire multiplier_0_n_32_110;
	 wire multiplier_0_n_32_111;
	 wire multiplier_0_n_32_112;
	 wire multiplier_0_n_32_113;
	 wire multiplier_0_n_32_114;
	 wire multiplier_0_n_32_115;
	 wire multiplier_0_n_32_116;
	 wire multiplier_0_n_32_117;
	 wire multiplier_0_n_32_118;
	 wire multiplier_0_n_32_119;
	 wire multiplier_0_n_32_120;
	 wire multiplier_0_n_32_121;
	 wire multiplier_0_n_32_122;
	 wire multiplier_0_n_32_123;
	 wire multiplier_0_n_32_124;
	 wire multiplier_0_n_32_125;
	 wire multiplier_0_n_32_126;
	 wire multiplier_0_n_32_127;
	 wire multiplier_0_n_32_128;
	 wire multiplier_0_n_32_129;
	 wire multiplier_0_n_32_130;
	 wire multiplier_0_n_32_131;
	 wire multiplier_0_n_32_132;
	 wire multiplier_0_n_32_133;
	 wire multiplier_0_n_32_134;
	 wire multiplier_0_n_32_135;
	 wire multiplier_0_n_32_136;
	 wire multiplier_0_n_32_137;
	 wire multiplier_0_n_32_138;
	 wire multiplier_0_n_32_139;
	 wire multiplier_0_n_32_140;
	 wire multiplier_0_n_32_141;
	 wire multiplier_0_n_32_142;
	 wire multiplier_0_n_32_143;
	 wire multiplier_0_n_32_144;
	 wire multiplier_0_n_32_145;
	 wire multiplier_0_n_32_146;
	 wire multiplier_0_n_32_147;
	 wire multiplier_0_n_32_148;
	 wire multiplier_0_n_32_149;
	 wire multiplier_0_n_32_150;
	 wire multiplier_0_n_32_151;
	 wire multiplier_0_n_32_152;
	 wire multiplier_0_n_32_153;
	 wire multiplier_0_n_32_154;
	 wire multiplier_0_n_32_155;
	 wire multiplier_0_n_32_156;
	 wire multiplier_0_n_32_157;
	 wire multiplier_0_n_32_158;
	 wire multiplier_0_n_32_159;
	 wire multiplier_0_n_32_160;
	 wire multiplier_0_n_32_161;
	 wire multiplier_0_n_32_162;
	 wire multiplier_0_n_32_163;
	 wire multiplier_0_n_32_164;
	 wire multiplier_0_n_32_165;
	 wire multiplier_0_n_32_166;
	 wire multiplier_0_n_32_167;
	 wire multiplier_0_n_32_168;
	 wire multiplier_0_n_32_169;
	 wire multiplier_0_n_32_170;
	 wire multiplier_0_n_32_171;
	 wire multiplier_0_n_32_172;
	 wire multiplier_0_n_32_173;
	 wire multiplier_0_n_32_174;
	 wire multiplier_0_n_32_175;
	 wire multiplier_0_n_32_176;
	 wire multiplier_0_n_32_177;
	 wire multiplier_0_n_32_178;
	 wire multiplier_0_n_32_179;
	 wire multiplier_0_n_32_180;
	 wire multiplier_0_n_32_181;
	 wire multiplier_0_n_32_182;
	 wire multiplier_0_n_32_183;
	 wire multiplier_0_n_32_184;
	 wire multiplier_0_n_32_185;
	 wire multiplier_0_n_32_186;
	 wire multiplier_0_n_32_187;
	 wire multiplier_0_n_32_188;
	 wire multiplier_0_n_32_189;
	 wire multiplier_0_n_32_190;
	 wire multiplier_0_n_32_191;
	 wire multiplier_0_n_32_192;
	 wire multiplier_0_n_32_193;
	 wire multiplier_0_n_32_194;
	 wire multiplier_0_n_32_195;
	 wire multiplier_0_n_32_196;
	 wire multiplier_0_n_32_197;
	 wire multiplier_0_n_32_198;
	 wire multiplier_0_n_32_199;
	 wire multiplier_0_n_32_200;
	 wire multiplier_0_n_32_201;
	 wire multiplier_0_n_32_202;
	 wire multiplier_0_n_32_203;
	 wire multiplier_0_n_32_204;
	 wire multiplier_0_n_32_205;
	 wire multiplier_0_n_32_206;
	 wire multiplier_0_n_32_207;
	 wire multiplier_0_n_32_208;
	 wire multiplier_0_n_32_209;
	 wire multiplier_0_n_32_210;
	 wire multiplier_0_n_32_211;
	 wire multiplier_0_n_32_212;
	 wire multiplier_0_n_32_213;
	 wire multiplier_0_n_32_214;
	 wire multiplier_0_n_32_215;
	 wire multiplier_0_n_32_216;
	 wire multiplier_0_n_32_217;
	 wire multiplier_0_n_32_218;
	 wire multiplier_0_n_32_219;
	 wire multiplier_0_n_32_220;
	 wire multiplier_0_n_32_221;
	 wire multiplier_0_n_32_222;
	 wire multiplier_0_n_32_223;
	 wire multiplier_0_n_32_224;
	 wire multiplier_0_n_32_225;
	 wire multiplier_0_n_32_226;
	 wire multiplier_0_n_32_227;
	 wire multiplier_0_n_32_228;
	 wire multiplier_0_n_32_229;
	 wire multiplier_0_n_32_230;
	 wire multiplier_0_n_32_231;
	 wire multiplier_0_n_32_232;
	 wire multiplier_0_n_32_233;
	 wire multiplier_0_n_32_234;
	 wire multiplier_0_n_32_235;
	 wire multiplier_0_n_32_236;
	 wire multiplier_0_n_32_237;
	 wire multiplier_0_n_32_238;
	 wire multiplier_0_n_32_239;
	 wire multiplier_0_n_32_240;
	 wire multiplier_0_n_32_241;
	 wire multiplier_0_n_32_242;
	 wire multiplier_0_n_32_243;
	 wire multiplier_0_n_32_244;
	 wire multiplier_0_n_32_245;
	 wire multiplier_0_n_32_246;
	 wire multiplier_0_n_32_247;
	 wire multiplier_0_n_32_248;
	 wire multiplier_0_n_32_249;
	 wire multiplier_0_n_32_250;
	 wire multiplier_0_n_32_251;
	 wire multiplier_0_n_32_252;
	 wire multiplier_0_n_32_253;
	 wire multiplier_0_n_32_254;
	 wire multiplier_0_n_32_255;
	 wire multiplier_0_n_32_256;
	 wire multiplier_0_n_32_257;
	 wire multiplier_0_n_32_258;
	 wire multiplier_0_n_32_259;
	 wire multiplier_0_n_32_260;
	 wire multiplier_0_n_32_261;
	 wire multiplier_0_n_32_262;
	 wire multiplier_0_n_32_263;
	 wire multiplier_0_n_32_264;
	 wire multiplier_0_n_32_265;
	 wire multiplier_0_n_32_266;
	 wire multiplier_0_n_32_267;
	 wire multiplier_0_n_32_268;
	 wire multiplier_0_n_32_269;
	 wire multiplier_0_n_32_270;
	 wire multiplier_0_n_32_271;
	 wire multiplier_0_n_32_272;
	 wire multiplier_0_n_32_273;
	 wire multiplier_0_n_32_274;
	 wire multiplier_0_n_32_275;
	 wire multiplier_0_n_32_276;
	 wire multiplier_0_n_32_277;
	 wire multiplier_0_n_32_278;
	 wire multiplier_0_n_32_279;
	 wire multiplier_0_n_32_280;
	 wire multiplier_0_n_32_281;
	 wire multiplier_0_n_32_282;
	 wire multiplier_0_n_32_283;
	 wire multiplier_0_n_32_284;
	 wire multiplier_0_n_32_285;
	 wire multiplier_0_n_32_286;
	 wire multiplier_0_n_32_287;
	 wire multiplier_0_n_32_288;
	 wire multiplier_0_n_32_289;
	 wire multiplier_0_n_32_290;
	 wire multiplier_0_n_32_291;
	 wire multiplier_0_n_32_292;
	 wire multiplier_0_n_32_293;
	 wire multiplier_0_n_32_294;
	 wire multiplier_0_n_32_295;
	 wire multiplier_0_n_32_296;
	 wire multiplier_0_n_32_297;
	 wire multiplier_0_n_32_298;
	 wire multiplier_0_n_32_299;
	 wire multiplier_0_n_32_300;
	 wire multiplier_0_n_32_301;
	 wire multiplier_0_n_32_302;
	 wire multiplier_0_n_32_303;
	 wire multiplier_0_n_32_304;
	 wire multiplier_0_n_32_305;
	 wire multiplier_0_n_32_306;
	 wire multiplier_0_n_32_307;
	 wire multiplier_0_n_32_308;
	 wire multiplier_0_n_32_309;
	 wire multiplier_0_n_32_310;
	 wire multiplier_0_n_32_311;
	 wire multiplier_0_n_32_312;
	 wire multiplier_0_n_32_313;
	 wire multiplier_0_n_32_314;
	 wire multiplier_0_n_32_315;
	 wire multiplier_0_n_32_316;
	 wire multiplier_0_n_32_317;
	 wire multiplier_0_n_32_318;
	 wire multiplier_0_n_32_319;
	 wire multiplier_0_n_32_320;
	 wire multiplier_0_n_32_321;
	 wire multiplier_0_n_32_322;
	 wire multiplier_0_n_32_323;
	 wire multiplier_0_n_32_324;
	 wire multiplier_0_n_32_325;
	 wire multiplier_0_n_32_326;
	 wire multiplier_0_n_32_327;
	 wire multiplier_0_n_32_328;
	 wire multiplier_0_n_32_329;
	 wire multiplier_0_n_32_330;
	 wire multiplier_0_n_32_331;
	 wire multiplier_0_n_32_332;
	 wire multiplier_0_n_32_333;
	 wire multiplier_0_n_32_334;
	 wire multiplier_0_n_32_335;
	 wire multiplier_0_n_32_336;
	 wire multiplier_0_n_32_337;
	 wire multiplier_0_n_32_338;
	 wire multiplier_0_n_32_339;
	 wire multiplier_0_n_32_340;
	 wire multiplier_0_n_32_341;
	 wire multiplier_0_n_32_342;
	 wire multiplier_0_n_32_343;
	 wire multiplier_0_n_32_344;
	 wire multiplier_0_n_32_345;
	 wire multiplier_0_n_32_346;
	 wire multiplier_0_n_32_347;
	 wire multiplier_0_n_32_348;
	 wire multiplier_0_n_32_349;
	 wire multiplier_0_n_32_350;
	 wire multiplier_0_n_32_351;
	 wire multiplier_0_n_32_352;
	 wire multiplier_0_n_32_353;
	 wire multiplier_0_n_32_354;
	 wire multiplier_0_n_32_355;
	 wire multiplier_0_n_32_356;
	 wire multiplier_0_n_32_357;
	 wire multiplier_0_n_32_358;
	 wire multiplier_0_n_32_359;
	 wire multiplier_0_n_32_360;
	 wire multiplier_0_n_32_361;
	 wire multiplier_0_n_32_362;
	 wire multiplier_0_n_32_363;
	 wire multiplier_0_n_32_364;
	 wire multiplier_0_n_32_365;
	 wire multiplier_0_n_32_366;
	 wire multiplier_0_n_32_367;
	 wire multiplier_0_n_32_368;
	 wire multiplier_0_n_32_369;
	 wire multiplier_0_n_32_370;
	 wire multiplier_0_n_32_371;
	 wire multiplier_0_n_32_372;
	 wire multiplier_0_n_32_373;
	 wire multiplier_0_n_32_374;
	 wire multiplier_0_n_32_375;
	 wire multiplier_0_n_32_376;
	 wire multiplier_0_n_32_377;
	 wire multiplier_0_n_32_378;
	 wire multiplier_0_n_32_379;
	 wire multiplier_0_n_32_380;
	 wire multiplier_0_n_32_381;
	 wire multiplier_0_n_32_382;
	 wire multiplier_0_n_32_383;
	 wire multiplier_0_n_32_384;
	 wire multiplier_0_n_32_385;
	 wire multiplier_0_n_32_386;
	 wire multiplier_0_n_32_387;
	 wire multiplier_0_n_32_388;
	 wire multiplier_0_n_32_389;
	 wire multiplier_0_n_32_390;
	 wire multiplier_0_n_32_391;
	 wire multiplier_0_n_32_392;
	 wire multiplier_0_n_32_393;
	 wire multiplier_0_n_32_394;
	 wire multiplier_0_n_32_395;
	 wire multiplier_0_n_32_396;
	 wire multiplier_0_n_32_397;
	 wire multiplier_0_n_32_398;
	 wire multiplier_0_n_32_399;
	 wire multiplier_0_n_32_400;
	 wire multiplier_0_n_32_401;
	 wire multiplier_0_n_32_402;
	 wire multiplier_0_n_32_403;
	 wire multiplier_0_n_32_404;
	 wire multiplier_0_n_32_405;
	 wire multiplier_0_n_32_406;
	 wire multiplier_0_n_32_407;
	 wire multiplier_0_n_32_408;
	 wire multiplier_0_n_32_409;
	 wire multiplier_0_n_32_410;
	 wire multiplier_0_n_32_411;
	 wire multiplier_0_n_32_412;
	 wire multiplier_0_n_32_413;
	 wire multiplier_0_n_32_414;
	 wire multiplier_0_n_32_415;
	 wire multiplier_0_n_32_416;
	 wire multiplier_0_n_32_417;
	 wire multiplier_0_n_32_418;
	 wire multiplier_0_n_32_419;
	 wire multiplier_0_n_32_420;
	 wire multiplier_0_n_32_421;
	 wire multiplier_0_n_32_422;
	 wire multiplier_0_n_32_423;
	 wire multiplier_0_n_32_424;
	 wire multiplier_0_n_32_425;
	 wire multiplier_0_n_32_426;
	 wire multiplier_0_n_32_427;
	 wire multiplier_0_n_32_428;
	 wire multiplier_0_n_32_429;
	 wire multiplier_0_n_32_430;
	 wire multiplier_0_n_32_431;
	 wire multiplier_0_n_32_432;
	 wire multiplier_0_n_32_433;
	 wire multiplier_0_n_32_434;
	 wire multiplier_0_n_32_435;
	 wire multiplier_0_n_32_436;
	 wire multiplier_0_n_32_437;
	 wire multiplier_0_n_32_438;
	 wire multiplier_0_n_32_439;
	 wire multiplier_0_n_32_440;
	 wire multiplier_0_n_32_441;
	 wire multiplier_0_n_32_442;
	 wire multiplier_0_n_32_443;
	 wire multiplier_0_n_32_444;
	 wire multiplier_0_n_32_445;
	 wire multiplier_0_n_32_446;
	 wire multiplier_0_n_32_447;
	 wire multiplier_0_n_32_448;
	 wire multiplier_0_n_32_449;
	 wire multiplier_0_n_32_450;
	 wire multiplier_0_n_32_451;
	 wire multiplier_0_n_32_452;
	 wire multiplier_0_n_32_453;
	 wire multiplier_0_n_32_454;
	 wire multiplier_0_n_32_455;
	 wire multiplier_0_n_32_456;
	 wire multiplier_0_n_32_457;
	 wire multiplier_0_n_32_458;
	 wire multiplier_0_n_32_459;
	 wire multiplier_0_n_32_460;
	 wire multiplier_0_n_32_461;
	 wire multiplier_0_n_32_462;
	 wire multiplier_0_n_32_463;
	 wire multiplier_0_n_32_464;
	 wire multiplier_0_n_32_465;
	 wire multiplier_0_n_32_466;
	 wire multiplier_0_n_32_467;
	 wire multiplier_0_n_32_468;
	 wire multiplier_0_n_32_469;
	 wire multiplier_0_n_32_470;
	 wire multiplier_0_n_32_471;
	 wire multiplier_0_n_32_472;
	 wire multiplier_0_n_32_473;
	 wire multiplier_0_n_32_474;
	 wire multiplier_0_n_32_475;
	 wire multiplier_0_n_32_476;
	 wire multiplier_0_n_32_477;
	 wire multiplier_0_n_32_478;
	 wire multiplier_0_n_32_479;
	 wire multiplier_0_n_32_480;
	 wire multiplier_0_n_32_481;
	 wire multiplier_0_n_32_482;
	 wire multiplier_0_n_32_483;
	 wire multiplier_0_n_32_484;
	 wire multiplier_0_n_32_485;
	 wire multiplier_0_n_32_486;
	 wire multiplier_0_n_32_487;
	 wire multiplier_0_n_32_488;
	 wire multiplier_0_n_32_489;
	 wire multiplier_0_n_32_490;
	 wire multiplier_0_n_32_491;
	 wire multiplier_0_n_32_492;
	 wire multiplier_0_n_32_493;
	 wire multiplier_0_n_32_494;
	 wire multiplier_0_n_32_495;
	 wire multiplier_0_n_32_496;
	 wire multiplier_0_n_32_497;
	 wire multiplier_0_n_32_498;
	 wire multiplier_0_n_32_499;
	 wire multiplier_0_n_32_500;
	 wire multiplier_0_n_32_501;
	 wire multiplier_0_n_32_502;
	 wire multiplier_0_n_32_503;
	 wire multiplier_0_n_32_504;
	 wire multiplier_0_n_32_505;
	 wire multiplier_0_n_32_506;
	 wire multiplier_0_n_32_507;
	 wire multiplier_0_n_32_508;
	 wire multiplier_0_n_32_509;
	 wire multiplier_0_n_32_510;
	 wire multiplier_0_n_32_511;
	 wire multiplier_0_n_32_512;
	 wire multiplier_0_n_32_513;
	 wire multiplier_0_n_32_514;
	 wire multiplier_0_n_32_515;
	 wire multiplier_0_n_32_516;
	 wire multiplier_0_n_32_517;
	 wire multiplier_0_n_32_518;
	 wire multiplier_0_n_32_519;
	 wire multiplier_0_n_32_520;
	 wire multiplier_0_n_32_521;
	 wire multiplier_0_n_32_522;
	 wire multiplier_0_n_32_523;
	 wire multiplier_0_n_32_524;
	 wire multiplier_0_n_32_525;
	 wire multiplier_0_n_32_526;
	 wire multiplier_0_n_32_527;
	 wire multiplier_0_n_32_528;
	 wire multiplier_0_n_32_529;
	 wire multiplier_0_n_32_530;
	 wire multiplier_0_n_32_531;
	 wire multiplier_0_n_32_532;
	 wire multiplier_0_n_32_533;
	 wire multiplier_0_n_32_534;
	 wire multiplier_0_n_32_535;
	 wire multiplier_0_n_32_536;
	 wire multiplier_0_n_32_537;
	 wire multiplier_0_n_32_538;
	 wire multiplier_0_n_32_539;
	 wire multiplier_0_n_32_540;
	 wire multiplier_0_n_32_541;
	 wire multiplier_0_n_32_542;
	 wire multiplier_0_n_32_543;
	 wire multiplier_0_n_32_544;
	 wire multiplier_0_n_32_545;
	 wire multiplier_0_n_32_546;
	 wire multiplier_0_n_32_547;
	 wire multiplier_0_n_32_548;
	 wire multiplier_0_n_32_549;
	 wire multiplier_0_n_32_550;
	 wire multiplier_0_n_32_551;
	 wire multiplier_0_n_32_552;
	 wire multiplier_0_n_32_553;
	 wire multiplier_0_n_32_554;
	 wire multiplier_0_n_32_555;
	 wire multiplier_0_n_32_556;
	 wire multiplier_0_n_32_557;
	 wire multiplier_0_n_32_558;
	 wire multiplier_0_n_32_559;
	 wire multiplier_0_n_32_560;
	 wire multiplier_0_n_32_561;
	 wire multiplier_0_n_32_562;
	 wire multiplier_0_n_32_563;
	 wire multiplier_0_n_32_564;
	 wire multiplier_0_n_32_565;
	 wire multiplier_0_n_32_566;
	 wire multiplier_0_n_32_567;
	 wire multiplier_0_n_32_568;
	 wire multiplier_0_n_32_569;
	 wire multiplier_0_n_32_570;
	 wire multiplier_0_n_32_571;
	 wire multiplier_0_n_32_572;
	 wire multiplier_0_n_32_573;
	 wire multiplier_0_n_32_574;
	 wire multiplier_0_n_32_575;
	 wire multiplier_0_n_32_576;
	 wire multiplier_0_n_32_577;
	 wire multiplier_0_n_32_578;
	 wire multiplier_0_n_32_579;
	 wire multiplier_0_n_32_580;
	 wire multiplier_0_n_32_581;
	 wire multiplier_0_n_32_582;
	 wire multiplier_0_n_32_583;
	 wire multiplier_0_n_32_584;
	 wire multiplier_0_n_32_585;
	 wire multiplier_0_n_32_586;
	 wire multiplier_0_n_32_587;
	 wire multiplier_0_n_32_588;
	 wire multiplier_0_n_32_589;
	 wire multiplier_0_n_32_590;
	 wire multiplier_0_n_32_591;
	 wire multiplier_0_n_32_592;
	 wire multiplier_0_n_32_593;
	 wire multiplier_0_n_32_594;
	 wire multiplier_0_n_32_595;
	 wire multiplier_0_n_32_596;
	 wire multiplier_0_n_32_597;
	 wire multiplier_0_n_32_598;
	 wire multiplier_0_n_32_599;
	 wire multiplier_0_n_32_600;
	 wire multiplier_0_n_32_601;
	 wire multiplier_0_n_32_602;
	 wire multiplier_0_n_32_603;
	 wire multiplier_0_n_32_604;
	 wire multiplier_0_n_32_605;
	 wire multiplier_0_n_32_606;
	 wire multiplier_0_n_32_607;
	 wire multiplier_0_n_32_608;
	 wire multiplier_0_n_32_609;
	 wire multiplier_0_n_32_610;
	 wire multiplier_0_n_32_611;
	 wire multiplier_0_n_32_612;
	 wire multiplier_0_n_32_613;
	 wire multiplier_0_n_32_614;
	 wire multiplier_0_n_32_615;
	 wire multiplier_0_n_32_616;
	 wire multiplier_0_n_32_617;
	 wire multiplier_0_n_32_618;
	 wire multiplier_0_n_32_619;
	 wire multiplier_0_n_32_620;
	 wire multiplier_0_n_32_621;
	 wire multiplier_0_n_32_622;
	 wire multiplier_0_n_32_623;
	 wire multiplier_0_n_32_624;
	 wire multiplier_0_n_32_625;
	 wire multiplier_0_n_32_626;
	 wire multiplier_0_n_32_627;
	 wire multiplier_0_n_32_628;
	 wire multiplier_0_n_32_629;
	 wire multiplier_0_n_32_630;
	 wire multiplier_0_n_32_631;
	 wire multiplier_0_n_32_632;
	 wire multiplier_0_n_32_633;
	 wire multiplier_0_n_32_634;
	 wire multiplier_0_n_32_635;
	 wire multiplier_0_n_32_636;
	 wire multiplier_0_n_32_637;
	 wire multiplier_0_n_32_638;
	 wire multiplier_0_n_32_639;
	 wire multiplier_0_n_32_640;
	 wire multiplier_0_n_32_641;
	 wire multiplier_0_n_32_642;
	 wire multiplier_0_n_32_643;
	 wire multiplier_0_n_32_644;
	 wire multiplier_0_n_32_645;
	 wire multiplier_0_n_32_646;
	 wire multiplier_0_n_32_647;
	 wire multiplier_0_n_32_648;
	 wire multiplier_0_n_32_649;
	 wire multiplier_0_n_32_650;
	 wire multiplier_0_n_32_651;
	 wire multiplier_0_n_32_652;
	 wire multiplier_0_n_32_653;
	 wire multiplier_0_n_32_654;
	 wire multiplier_0_n_32_655;
	 wire multiplier_0_n_32_656;
	 wire multiplier_0_n_32_657;
	 wire multiplier_0_n_32_658;
	 wire multiplier_0_n_32_659;
	 wire multiplier_0_n_32_660;
	 wire multiplier_0_n_32_661;
	 wire multiplier_0_n_32_662;
	 wire multiplier_0_n_32_663;
	 wire multiplier_0_n_32_664;
	 wire multiplier_0_n_32_665;
	 wire multiplier_0_n_32_666;
	 wire multiplier_0_n_32_667;
	 wire multiplier_0_n_32_668;
	 wire multiplier_0_n_32_669;
	 wire multiplier_0_n_32_670;
	 wire multiplier_0_n_32_671;
	 wire multiplier_0_n_32_672;
	 wire multiplier_0_n_32_673;
	 wire multiplier_0_n_32_674;
	 wire multiplier_0_n_34_0;
	 wire [31:0]multiplier_0_product_xp;
	 wire multiplier_0_n_34_1;
	 wire multiplier_0_n_34_2;
	 wire multiplier_0_n_34_3;
	 wire multiplier_0_n_34_4;
	 wire multiplier_0_n_34_5;
	 wire multiplier_0_n_34_6;
	 wire multiplier_0_n_34_7;
	 wire multiplier_0_n_34_8;
	 wire multiplier_0_n_34_9;
	 wire multiplier_0_n_34_10;
	 wire multiplier_0_n_34_11;
	 wire multiplier_0_n_34_12;
	 wire multiplier_0_n_34_13;
	 wire multiplier_0_n_34_14;
	 wire multiplier_0_n_34_15;
	 wire multiplier_0_n_34_16;
	 wire multiplier_0_n_34_17;
	 wire multiplier_0_n_34_18;
	 wire multiplier_0_n_34_19;
	 wire multiplier_0_n_34_20;
	 wire multiplier_0_n_34_21;
	 wire multiplier_0_n_34_22;
	 wire multiplier_0_n_34_23;
	 wire multiplier_0_n_34_24;
	 wire multiplier_0_n_34_25;
	 wire multiplier_0_acc_sel;
	 wire multiplier_0_n_38_0;
	 wire multiplier_0_result_clr;
	 wire multiplier_0_n_39_0;
	 wire multiplier_0_n_39_1;
	 wire [15:0]multiplier_0_reshi;
	 wire multiplier_0_n_41_0;
	 wire multiplier_0_n_41_1;
	 wire multiplier_0_n_41_2;
	 wire multiplier_0_n_41_3;
	 wire multiplier_0_n_41_4;
	 wire multiplier_0_n_41_5;
	 wire multiplier_0_n_41_6;
	 wire multiplier_0_n_41_7;
	 wire multiplier_0_n_41_8;
	 wire multiplier_0_n_41_9;
	 wire multiplier_0_n_41_10;
	 wire multiplier_0_n_41_11;
	 wire multiplier_0_n_41_12;
	 wire multiplier_0_n_41_13;
	 wire multiplier_0_n_41_14;
	 wire multiplier_0_n_41_15;
	 wire multiplier_0_n_41_16;
	 wire multiplier_0_n_42_0;
	 wire multiplier_0_n_42_1;
	 wire multiplier_0_n_45_0;
	 wire multiplier_0_n_45_1;
	 wire multiplier_0_n_45_2;
	 wire multiplier_0_n_45_3;
	 wire multiplier_0_n_45_4;
	 wire multiplier_0_n_45_5;
	 wire multiplier_0_n_45_6;
	 wire multiplier_0_n_45_7;
	 wire multiplier_0_n_45_8;
	 wire multiplier_0_n_45_9;
	 wire multiplier_0_n_45_10;
	 wire multiplier_0_n_45_11;
	 wire multiplier_0_n_45_12;
	 wire multiplier_0_n_45_13;
	 wire multiplier_0_n_45_14;
	 wire multiplier_0_n_45_15;
	 wire multiplier_0_n_45_16;
	 wire multiplier_0_n_46_0;
	 wire multiplier_0_n_46_1;
	 wire multiplier_0_n_48_0;
	 wire multiplier_0_n_48_1;
	 wire multiplier_0_n_48_2;
	 wire multiplier_0_n_48_3;
	 wire multiplier_0_n_48_4;
	 wire multiplier_0_n_48_5;
	 wire multiplier_0_n_48_6;
	 wire multiplier_0_n_48_7;
	 wire multiplier_0_n_48_8;
	 wire multiplier_0_n_48_9;
	 wire multiplier_0_n_48_10;
	 wire multiplier_0_n_48_11;
	 wire multiplier_0_n_48_12;
	 wire multiplier_0_n_48_13;
	 wire multiplier_0_n_48_14;
	 wire multiplier_0_n_48_15;
	 wire [15:0]multiplier_0_reshi_nxt;
	 wire multiplier_0_n_48_16;
	 wire multiplier_0_n_48_17;
	 wire multiplier_0_n_48_18;
	 wire multiplier_0_n_48_19;
	 wire multiplier_0_n_48_20;
	 wire multiplier_0_n_48_21;
	 wire multiplier_0_n_48_22;
	 wire multiplier_0_n_48_23;
	 wire multiplier_0_n_48_24;
	 wire multiplier_0_n_48_25;
	 wire multiplier_0_n_48_26;
	 wire multiplier_0_n_48_27;
	 wire multiplier_0_n_48_28;
	 wire multiplier_0_n_48_29;
	 wire multiplier_0_n_48_30;
	 wire multiplier_0_n_50_0;
	 wire multiplier_0_n_50_1;
	 wire [1:0]multiplier_0_sumext_s_nxt;
	 wire [1:0]multiplier_0_sumext_s;
	 wire multiplier_0_n_52_0;
	 wire multiplier_0_n_53_0;
	 wire multiplier_0_n_53_1;
	 wire multiplier_0_n_55_0;
	 wire multiplier_0_n_55_1;
	 wire multiplier_0_n_55_2;
	 wire multiplier_0_n_57_0;
	 wire multiplier_0_n_57_1;
	 wire multiplier_0_n_60_0;
	 wire multiplier_0_n_60_1;
	 wire multiplier_0_n_60_2;
	 wire multiplier_0_n_60_3;
	 wire multiplier_0_n_60_4;
	 wire multiplier_0_n_60_5;
	 wire multiplier_0_n_60_6;
	 wire multiplier_0_n_60_7;
	 wire multiplier_0_n_60_8;
	 wire multiplier_0_n_60_9;
	 wire multiplier_0_n_60_10;
	 wire multiplier_0_n_60_11;
	 wire multiplier_0_n_60_12;
	 wire multiplier_0_n_60_13;
	 wire multiplier_0_n_60_14;
	 wire multiplier_0_n_60_15;
	 wire multiplier_0_n_60_16;
	 wire multiplier_0_n_60_17;
	 wire multiplier_0_n_60_18;
	 wire multiplier_0_n_60_19;
	 wire multiplier_0_n_60_20;
	 wire multiplier_0_n_60_21;
	 wire multiplier_0_n_60_22;
	 wire multiplier_0_n_60_23;
	 wire multiplier_0_n_60_24;
	 wire multiplier_0_n_60_25;
	 wire multiplier_0_n_60_26;
	 wire multiplier_0_n_60_27;
	 wire multiplier_0_n_60_28;
	 wire multiplier_0_n_60_29;
	 wire multiplier_0_n_60_30;
	 wire multiplier_0_n_60_31;
	 wire multiplier_0_n_60_32;
	 wire multiplier_0_n_60_33;
	 wire multiplier_0_n_60_34;
	 wire multiplier_0_n_60_35;
	 wire multiplier_0_n_60_36;
	 wire multiplier_0_n_60_37;
	 wire multiplier_0_n_60_38;
	 wire multiplier_0_n_60_39;
	 wire multiplier_0_n_60_40;
	 wire multiplier_0_n_60_41;
	 wire multiplier_0_n_60_42;
	 wire multiplier_0_n_60_43;
	 wire multiplier_0_n_60_44;
	 wire multiplier_0_n_60_45;
	 wire multiplier_0_n_60_46;
	 wire multiplier_0_n_60_47;
	 wire multiplier_0_n_60_48;
	 wire multiplier_0_n_60_49;
	 wire multiplier_0_n_60_50;
	 wire multiplier_0_n_60_51;
	 wire multiplier_0_n_60_52;
	 wire multiplier_0_n_60_53;
	 wire multiplier_0_n_60_54;
	 wire multiplier_0_n_60_55;
	 wire multiplier_0_n_60_56;
	 wire multiplier_0_n_60_57;
	 wire multiplier_0_n_60_58;
	 wire multiplier_0_n_60_59;
	 wire multiplier_0_n_60_60;
	 wire multiplier_0_n_60_61;
	 wire multiplier_0_n_60_62;
	 wire multiplier_0_n_60_63;
	 wire multiplier_0_n_60_64;
	 wire multiplier_0_n_60_65;
	 wire multiplier_0_n_60_66;
	 wire multiplier_0_n_60_67;
	 wire multiplier_0_n_60_68;
	 wire multiplier_0_n_60_69;
	 wire multiplier_0_n_60_70;
	 wire multiplier_0_n_60_71;
	 wire multiplier_0_n_60_72;
	 wire multiplier_0_n_60_73;
	 wire multiplier_0_n_60_74;
	 wire multiplier_0_n_60_75;
	 wire multiplier_0_n_60_76;
	 wire multiplier_0_n_60_77;
	 wire multiplier_0_n_60_78;
	 wire multiplier_0_n_60_79;
	 wire multiplier_0_n_60_80;
	 wire multiplier_0_n_60_81;
	 wire multiplier_0_n_60_82;
	 wire multiplier_0_n_15;
	 wire multiplier_0_n_5;
	 wire multiplier_0_n_38;
	 wire multiplier_0_n_3;
	 wire multiplier_0_n_18;
	 wire multiplier_0_n_4;
	 wire multiplier_0_n_19;
	 wire multiplier_0_n_68;
	 wire multiplier_0_n_1;
	 wire multiplier_0_n_16;
	 wire multiplier_0_n_2;
	 wire multiplier_0_n_17;
	 wire multiplier_0_n_67;
	 wire multiplier_0_n_6;
	 wire multiplier_0_n_20;
	 wire multiplier_0_n_21;
	 wire multiplier_0_n_41;
	 wire multiplier_0_n_45;
	 wire multiplier_0_n_46;
	 wire multiplier_0_n_47;
	 wire multiplier_0_n_48;
	 wire multiplier_0_n_49;
	 wire multiplier_0_n_40;
	 wire multiplier_0_n_39;
	 wire multiplier_0_n_50;
	 wire multiplier_0_n_51;
	 wire multiplier_0_n_52;
	 wire multiplier_0_n_53;
	 wire multiplier_0_n_54;
	 wire multiplier_0_n_55;
	 wire multiplier_0_n_56;
	 wire multiplier_0_n_57;
	 wire multiplier_0_n_136;
	 wire multiplier_0_n_119;
	 wire multiplier_0_n_69;
	 wire multiplier_0_n_121;
	 wire multiplier_0_n_88;
	 wire multiplier_0_n_90;
	 wire multiplier_0_n_135;
	 wire multiplier_0_n_118;
	 wire multiplier_0_n_91;
	 wire multiplier_0_n_134;
	 wire multiplier_0_n_117;
	 wire multiplier_0_n_92;
	 wire multiplier_0_n_133;
	 wire multiplier_0_n_116;
	 wire multiplier_0_n_93;
	 wire multiplier_0_n_44;
	 wire multiplier_0_n_132;
	 wire multiplier_0_n_115;
	 wire multiplier_0_n_94;
	 wire multiplier_0_n_43;
	 wire multiplier_0_n_131;
	 wire multiplier_0_n_114;
	 wire multiplier_0_n_95;
	 wire multiplier_0_n_42;
	 wire multiplier_0_n_130;
	 wire multiplier_0_n_113;
	 wire multiplier_0_n_96;
	 wire multiplier_0_n_129;
	 wire multiplier_0_n_112;
	 wire multiplier_0_n_97;
	 wire multiplier_0_n_128;
	 wire multiplier_0_n_111;
	 wire multiplier_0_n_98;
	 wire multiplier_0_n_127;
	 wire multiplier_0_n_110;
	 wire multiplier_0_n_99;
	 wire multiplier_0_n_126;
	 wire multiplier_0_n_109;
	 wire multiplier_0_n_100;
	 wire multiplier_0_n_125;
	 wire multiplier_0_n_108;
	 wire multiplier_0_n_101;
	 wire multiplier_0_n_124;
	 wire multiplier_0_n_107;
	 wire multiplier_0_n_102;
	 wire multiplier_0_n_123;
	 wire multiplier_0_n_106;
	 wire multiplier_0_n_103;
	 wire multiplier_0_n_122;
	 wire multiplier_0_n_105;
	 wire multiplier_0_n_104;
	 wire multiplier_0_n_89;
	 wire multiplier_0_n_137;
	 wire multiplier_0_n_120;
	 wire multiplier_0_n_0;
	 wire multiplier_0_n_13;
	 wire multiplier_0_n_9;
	 wire multiplier_0_n_11;
	 wire multiplier_0_n_10;
	 wire multiplier_0_n_150;
	 wire multiplier_0_n_58;
	 wire multiplier_0_n_59;
	 wire multiplier_0_n_60;
	 wire multiplier_0_n_61;
	 wire multiplier_0_n_62;
	 wire multiplier_0_n_63;
	 wire multiplier_0_n_64;
	 wire multiplier_0_n_65;
	 wire multiplier_0_n_66;
	 wire multiplier_0_n_7;
	 wire multiplier_0_n_86;
	 wire multiplier_0_n_87;
	 wire multiplier_0_n_70;
	 wire multiplier_0_n_85;
	 wire multiplier_0_n_84;
	 wire multiplier_0_n_83;
	 wire multiplier_0_n_82;
	 wire multiplier_0_n_81;
	 wire multiplier_0_n_80;
	 wire multiplier_0_n_79;
	 wire multiplier_0_n_78;
	 wire multiplier_0_n_77;
	 wire multiplier_0_n_76;
	 wire multiplier_0_n_75;
	 wire multiplier_0_n_74;
	 wire multiplier_0_n_73;
	 wire multiplier_0_n_72;
	 wire multiplier_0_n_71;
	 wire multiplier_0_n_138;
	 wire multiplier_0_n_142;
	 wire multiplier_0_n_143;
	 wire multiplier_0_n_140;
	 wire multiplier_0_n_148;
	 wire multiplier_0_n_8;
	 wire multiplier_0_n_149;
	 wire multiplier_0_n_12;
	 wire multiplier_0_n_37;
	 wire multiplier_0_n_14;
	 wire multiplier_0_n_36;
	 wire multiplier_0_n_35;
	 wire multiplier_0_n_34;
	 wire multiplier_0_n_33;
	 wire multiplier_0_n_32;
	 wire multiplier_0_n_31;
	 wire multiplier_0_n_30;
	 wire multiplier_0_n_29;
	 wire multiplier_0_n_28;
	 wire multiplier_0_n_27;
	 wire multiplier_0_n_26;
	 wire multiplier_0_n_25;
	 wire multiplier_0_n_24;
	 wire multiplier_0_n_145;
	 wire multiplier_0_n_147;
	 wire multiplier_0_n_23;
	 wire multiplier_0_n_139;
	 wire multiplier_0_n_141;
	 wire multiplier_0_n_144;
	 wire multiplier_0_n_146;
	 wire multiplier_0_n_22;
	 wire mem_backbone_0_n_0_0;
	 wire [15:0]mem_backbone_0_per_dout_val;
	 wire mem_backbone_0_n_2_0;
	 wire mem_backbone_0_n_2_1;
	 wire [14:0]mem_backbone_0_ext_mem_addr;
	 wire mem_backbone_0_n_2_2;
	 wire mem_backbone_0_n_2_3;
	 wire mem_backbone_0_n_2_4;
	 wire mem_backbone_0_n_2_5;
	 wire mem_backbone_0_n_2_6;
	 wire mem_backbone_0_n_2_7;
	 wire mem_backbone_0_n_2_8;
	 wire mem_backbone_0_n_2_9;
	 wire mem_backbone_0_n_2_10;
	 wire mem_backbone_0_n_2_11;
	 wire mem_backbone_0_n_2_12;
	 wire mem_backbone_0_n_2_13;
	 wire mem_backbone_0_n_2_14;
	 wire mem_backbone_0_n_2_15;
	 wire mem_backbone_0_n_3_0;
	 wire mem_backbone_0_ext_per_sel;
	 wire mem_backbone_0_ext_mem_en;
	 wire mem_backbone_0_n_5_0;
	 wire mem_backbone_0_n_5_1;
	 wire mem_backbone_0_n_5_2;
	 wire mem_backbone_0_eu_per_en;
	 wire mem_backbone_0_n_6_0;
	 wire mem_backbone_0_ext_per_en;
	 wire mem_backbone_0_ext_pmem_sel;
	 wire mem_backbone_0_n_8_0;
	 wire mem_backbone_0_fe_pmem_en;
	 wire mem_backbone_0_n_11_0;
	 wire mem_backbone_0_n_11_1;
	 wire mem_backbone_0_eu_pmem_en;
	 wire mem_backbone_0_n_12_0;
	 wire mem_backbone_0_ext_pmem_en;
	 wire [1:0]mem_backbone_0_ext_mem_din_sel;
	 wire mem_backbone_0_n_15_0;
	 wire mem_backbone_0_n_16_0;
	 wire mem_backbone_0_n_16_1;
	 wire mem_backbone_0_n_16_2;
	 wire mem_backbone_0_n_16_3;
	 wire mem_backbone_0_n_16_4;
	 wire mem_backbone_0_n_16_5;
	 wire mem_backbone_0_n_16_6;
	 wire mem_backbone_0_n_16_7;
	 wire mem_backbone_0_n_16_8;
	 wire mem_backbone_0_n_16_9;
	 wire mem_backbone_0_n_16_10;
	 wire mem_backbone_0_n_16_11;
	 wire mem_backbone_0_n_16_12;
	 wire mem_backbone_0_n_16_13;
	 wire mem_backbone_0_n_16_14;
	 wire mem_backbone_0_n_16_15;
	 wire mem_backbone_0_n_19_0;
	 wire mem_backbone_0_n_19_1;
	 wire mem_backbone_0_n_19_2;
	 wire mem_backbone_0_n_19_3;
	 wire mem_backbone_0_n_19_4;
	 wire mem_backbone_0_n_19_5;
	 wire mem_backbone_0_n_19_6;
	 wire mem_backbone_0_ext_dmem_sel;
	 wire mem_backbone_0_n_20_0;
	 wire mem_backbone_0_n_20_1;
	 wire mem_backbone_0_n_20_2;
	 wire mem_backbone_0_n_20_3;
	 wire mem_backbone_0_n_20_4;
	 wire mem_backbone_0_n_20_5;
	 wire mem_backbone_0_eu_dmem_en;
	 wire mem_backbone_0_n_21_0;
	 wire mem_backbone_0_ext_dmem_en;
	 wire mem_backbone_0_n_22_0;
	 wire mem_backbone_0_n_22_1;
	 wire mem_backbone_0_n_22_2;
	 wire mem_backbone_0_n_22_3;
	 wire mem_backbone_0_n_22_4;
	 wire mem_backbone_0_n_22_5;
	 wire mem_backbone_0_n_22_6;
	 wire mem_backbone_0_n_22_7;
	 wire mem_backbone_0_n_22_8;
	 wire mem_backbone_0_n_22_9;
	 wire mem_backbone_0_n_24_0;
	 wire mem_backbone_0_n_24_1;
	 wire mem_backbone_0_n_24_2;
	 wire mem_backbone_0_n_24_3;
	 wire mem_backbone_0_n_24_4;
	 wire mem_backbone_0_n_24_5;
	 wire mem_backbone_0_n_24_6;
	 wire mem_backbone_0_n_24_7;
	 wire mem_backbone_0_n_24_8;
	 wire mem_backbone_0_n_24_9;
	 wire mem_backbone_0_n_24_10;
	 wire mem_backbone_0_n_24_11;
	 wire mem_backbone_0_n_24_12;
	 wire mem_backbone_0_n_24_13;
	 wire mem_backbone_0_n_24_14;
	 wire mem_backbone_0_n_24_15;
	 wire mem_backbone_0_n_24_16;
	 wire mem_backbone_0_n_25_0;
	 wire mem_backbone_0_n_25_1;
	 wire mem_backbone_0_n_25_2;
	 wire mem_backbone_0_n_25_3;
	 wire mem_backbone_0_n_25_4;
	 wire mem_backbone_0_n_25_5;
	 wire mem_backbone_0_n_25_6;
	 wire mem_backbone_0_n_25_7;
	 wire mem_backbone_0_n_25_8;
	 wire mem_backbone_0_n_25_9;
	 wire mem_backbone_0_n_25_10;
	 wire mem_backbone_0_n_25_11;
	 wire mem_backbone_0_n_25_12;
	 wire mem_backbone_0_n_25_13;
	 wire mem_backbone_0_n_25_14;
	 wire mem_backbone_0_n_25_15;
	 wire mem_backbone_0_n_25_16;
	 wire mem_backbone_0_n_27_0;
	 wire mem_backbone_0_n_27_1;
	 wire [1:0]mem_backbone_0_ext_mem_wr;
	 wire mem_backbone_0_n_27_2;
	 wire mem_backbone_0_n_29_0;
	 wire mem_backbone_0_n_29_1;
	 wire mem_backbone_0_n_29_2;
	 wire [1:0]mem_backbone_0_eu_mdb_in_sel;
	 wire mem_backbone_0_n_31_0;
	 wire mem_backbone_0_n_32_0;
	 wire mem_backbone_0_n_32_1;
	 wire mem_backbone_0_n_32_2;
	 wire mem_backbone_0_n_32_3;
	 wire mem_backbone_0_n_32_4;
	 wire mem_backbone_0_n_32_5;
	 wire mem_backbone_0_n_32_6;
	 wire mem_backbone_0_n_32_7;
	 wire mem_backbone_0_n_32_8;
	 wire mem_backbone_0_n_32_9;
	 wire mem_backbone_0_n_32_10;
	 wire mem_backbone_0_n_32_11;
	 wire mem_backbone_0_n_32_12;
	 wire mem_backbone_0_n_32_13;
	 wire mem_backbone_0_n_32_14;
	 wire mem_backbone_0_n_32_15;
	 wire mem_backbone_0_fe_pmem_en_dly;
	 wire mem_backbone_0_n_33_0;
	 wire mem_backbone_0_fe_pmem_save;
	 wire [15:0]mem_backbone_0_pmem_dout_bckup;
	 wire mem_backbone_0_n_35_0;
	 wire mem_backbone_0_n_35_1;
	 wire mem_backbone_0_fe_pmem_restore;
	 wire mem_backbone_0_pmem_dout_bckup_sel;
	 wire mem_backbone_0_n_37_0;
	 wire mem_backbone_0_n_37_1;
	 wire mem_backbone_0_n_39_0;
	 wire mem_backbone_0_n_39_1;
	 wire mem_backbone_0_n_39_2;
	 wire mem_backbone_0_n_39_3;
	 wire mem_backbone_0_n_39_4;
	 wire mem_backbone_0_n_39_5;
	 wire mem_backbone_0_n_39_6;
	 wire mem_backbone_0_n_39_7;
	 wire mem_backbone_0_n_39_8;
	 wire mem_backbone_0_n_39_9;
	 wire mem_backbone_0_n_39_10;
	 wire mem_backbone_0_n_39_11;
	 wire mem_backbone_0_n_39_12;
	 wire mem_backbone_0_n_39_13;
	 wire mem_backbone_0_n_39_14;
	 wire mem_backbone_0_n_39_15;
	 wire mem_backbone_0_n_39_16;
	 wire mem_backbone_0_n_42_0;
	 wire mem_backbone_0_n_43_0;
	 wire mem_backbone_0_dma_ready_dly;
	 wire mem_backbone_0_n_45_0;
	 wire mem_backbone_0_n_45_1;
	 wire mem_backbone_0_n_45_2;
	 wire mem_backbone_0_n_45_3;
	 wire mem_backbone_0_n_45_4;
	 wire mem_backbone_0_n_45_5;
	 wire mem_backbone_0_n_45_6;
	 wire mem_backbone_0_n_45_7;
	 wire mem_backbone_0_n_45_8;
	 wire mem_backbone_0_n_46_0;
	 wire mem_backbone_0_n_46_1;
	 wire mem_backbone_0_n_46_2;
	 wire mem_backbone_0_n_46_3;
	 wire mem_backbone_0_n_46_4;
	 wire mem_backbone_0_n_46_5;
	 wire mem_backbone_0_n_46_6;
	 wire mem_backbone_0_n_46_7;
	 wire mem_backbone_0_n_46_8;
	 wire mem_backbone_0_n_46_9;
	 wire mem_backbone_0_n_46_10;
	 wire mem_backbone_0_n_46_11;
	 wire mem_backbone_0_n_46_12;
	 wire mem_backbone_0_n_46_13;
	 wire mem_backbone_0_n_46_14;
	 wire mem_backbone_0_n_46_15;
	 wire mem_backbone_0_n_46_16;
	 wire mem_backbone_0_n_47_0;
	 wire mem_backbone_0_n_47_1;
	 wire mem_backbone_0_n_47_2;
	 wire mem_backbone_0_n_49_0;
	 wire mem_backbone_0_n_49_1;
	 wire mem_backbone_0_n_49_2;
	 wire mem_backbone_0_n_49_3;
	 wire mem_backbone_0_n_49_4;
	 wire mem_backbone_0_n_49_5;
	 wire mem_backbone_0_n_49_6;
	 wire mem_backbone_0_n_49_7;
	 wire mem_backbone_0_n_49_8;
	 wire mem_backbone_0_n_49_9;
	 wire mem_backbone_0_n_49_10;
	 wire mem_backbone_0_n_49_11;
	 wire mem_backbone_0_n_51_0;
	 wire mem_backbone_0_n_51_1;
	 wire mem_backbone_0_n_0;
	 wire mem_backbone_0_n_1;
	 wire mem_backbone_0_n_2;
	 wire mem_backbone_0_n_4;
	 wire mem_backbone_0_n_3;
	 wire mem_backbone_0_n_5;
	 wire mem_backbone_0_n_6;
	 wire mem_backbone_0_n_8;
	 wire mem_backbone_0_n_10;
	 wire mem_backbone_0_n_7;
	 wire mem_backbone_0_n_9;
	 wire mem_backbone_0_n_12;
	 wire mem_backbone_0_n_11;
	 wire mem_backbone_0_n_15;
	 wire mem_backbone_0_n_14;
	 wire mem_backbone_0_n_13;
	 wire mem_backbone_0_n_16;
	 wire frontend_0_mirq_wkup;
	 wire frontend_0_n_0_0;
	 wire frontend_0_cpu_halt_req;
	 wire frontend_0_n_3_0;
	 wire frontend_0_n_3_1;
	 wire frontend_0_n_3_2;
	 wire frontend_0_n_3_3;
	 wire frontend_0_n_4_0;
	 wire frontend_0_n_4_1;
	 wire frontend_0_n_4_2;
	 wire [2:0]frontend_0_i_state;
	 wire frontend_0_n_6_0;
	 wire frontend_0_n_6_1;
	 wire frontend_0_n_6_2;
	 wire frontend_0_n_10_0;
	 wire frontend_0_n_10_1;
	 wire [3:0]frontend_0_src_reg;
	 wire frontend_0_n_10_2;
	 wire frontend_0_n_10_3;
	 wire frontend_0_n_10_4;
	 wire frontend_0_n_11_0;
	 wire frontend_0_inst_type_nxt;
	 wire frontend_0_n_12_0;
	 wire frontend_0_n_12_1;
	 wire frontend_0_n_12_2;
	 wire frontend_0_n_12_3;
	 wire frontend_0_n_12_4;
	 wire frontend_0_n_12_5;
	 wire frontend_0_n_12_6;
	 wire frontend_0_n_12_7;
	 wire frontend_0_n_12_8;
	 wire frontend_0_n_12_9;
	 wire [12:0]frontend_0_inst_as_nxt;
	 wire frontend_0_n_12_10;
	 wire frontend_0_n_12_11;
	 wire frontend_0_n_12_12;
	 wire frontend_0_n_12_13;
	 wire frontend_0_n_12_14;
	 wire frontend_0_n_13_0;
	 wire frontend_0_n_13_1;
	 wire frontend_0_is_const;
	 wire frontend_0_is_sext;
	 wire frontend_0_n_16_0;
	 wire frontend_0_inst_dext_rdy;
	 wire frontend_0_exec_dext_rdy;
	 wire frontend_0_n_19_0;
	 wire frontend_0_n_19_1;
	 wire frontend_0_n_20_0;
	 wire frontend_0_n_20_1;
	 wire frontend_0_n_20_2;
	 wire frontend_0_n_20_3;
	 wire frontend_0_n_22_0;
	 wire frontend_0_n_23_0;
	 wire frontend_0_n_23_1;
	 wire frontend_0_n_23_2;
	 wire frontend_0_n_23_3;
	 wire frontend_0_n_23_4;
	 wire frontend_0_n_23_5;
	 wire frontend_0_n_23_6;
	 wire frontend_0_n_23_7;
	 wire frontend_0_n_23_8;
	 wire frontend_0_n_23_9;
	 wire frontend_0_n_23_10;
	 wire frontend_0_n_23_11;
	 wire frontend_0_n_23_12;
	 wire frontend_0_n_23_13;
	 wire frontend_0_n_23_14;
	 wire frontend_0_n_23_15;
	 wire frontend_0_n_23_16;
	 wire frontend_0_n_23_17;
	 wire frontend_0_inst_ad_nxt;
	 wire frontend_0_n_25_0;
	 wire frontend_0_n_25_1;
	 wire frontend_0_n_25_2;
	 wire frontend_0_n_25_3;
	 wire frontend_0_n_25_4;
	 wire frontend_0_n_25_5;
	 wire frontend_0_n_25_6;
	 wire frontend_0_n_27_0;
	 wire [7:0]frontend_0_inst_so_nxt;
	 wire frontend_0_n_27_1;
	 wire frontend_0_inst_sext_rdy;
	 wire frontend_0_exec_dst_wr;
	 wire frontend_0_n_32_0;
	 wire frontend_0_n_33_0;
	 wire frontend_0_n_33_1;
	 wire frontend_0_n_33_2;
	 wire frontend_0_n_33_3;
	 wire frontend_0_n_33_4;
	 wire frontend_0_exec_src_wr;
	 wire frontend_0_n_39_0;
	 wire frontend_0_n_39_1;
	 wire frontend_0_exec_jmp;
	 wire frontend_0_n_44_0;
	 wire frontend_0_n_44_1;
	 wire frontend_0_n_45_0;
	 wire frontend_0_n_45_1;
	 wire frontend_0_n_45_2;
	 wire frontend_0_dst_acalc_pre;
	 wire frontend_0_src_acalc_pre;
	 wire frontend_0_n_50_0;
	 wire frontend_0_n_50_1;
	 wire frontend_0_n_50_2;
	 wire frontend_0_n_50_3;
	 wire frontend_0_n_50_4;
	 wire frontend_0_n_50_5;
	 wire frontend_0_n_50_6;
	 wire frontend_0_n_50_7;
	 wire frontend_0_n_50_8;
	 wire frontend_0_n_50_9;
	 wire frontend_0_n_50_10;
	 wire frontend_0_n_50_11;
	 wire frontend_0_n_50_12;
	 wire frontend_0_n_50_13;
	 wire frontend_0_n_50_14;
	 wire frontend_0_n_50_15;
	 wire frontend_0_n_50_16;
	 wire frontend_0_n_50_17;
	 wire frontend_0_n_50_18;
	 wire frontend_0_n_50_19;
	 wire frontend_0_n_53_0;
	 wire frontend_0_n_53_1;
	 wire frontend_0_n_55_0;
	 wire frontend_0_n_55_1;
	 wire frontend_0_n_55_2;
	 wire frontend_0_n_55_3;
	 wire frontend_0_n_55_4;
	 wire frontend_0_n_55_5;
	 wire frontend_0_n_55_6;
	 wire frontend_0_n_55_7;
	 wire frontend_0_n_55_8;
	 wire frontend_0_n_55_9;
	 wire frontend_0_n_55_10;
	 wire frontend_0_n_55_11;
	 wire frontend_0_n_55_12;
	 wire frontend_0_n_55_13;
	 wire frontend_0_n_55_14;
	 wire frontend_0_n_55_15;
	 wire frontend_0_n_55_16;
	 wire frontend_0_n_55_17;
	 wire frontend_0_n_55_18;
	 wire frontend_0_n_55_19;
	 wire frontend_0_n_55_20;
	 wire frontend_0_n_55_21;
	 wire frontend_0_n_55_22;
	 wire frontend_0_n_55_23;
	 wire frontend_0_n_55_24;
	 wire frontend_0_n_55_25;
	 wire frontend_0_n_55_26;
	 wire frontend_0_n_55_27;
	 wire frontend_0_n_55_28;
	 wire frontend_0_n_55_29;
	 wire frontend_0_n_55_30;
	 wire frontend_0_n_55_31;
	 wire frontend_0_n_55_32;
	 wire frontend_0_n_55_33;
	 wire frontend_0_n_55_34;
	 wire [3:0]frontend_0_e_state_nxt_reg;
	 wire frontend_0_n_55_35;
	 wire frontend_0_n_55_36;
	 wire frontend_0_n_55_37;
	 wire frontend_0_n_55_38;
	 wire frontend_0_n_55_39;
	 wire frontend_0_n_55_40;
	 wire frontend_0_n_55_41;
	 wire frontend_0_n_55_42;
	 wire frontend_0_n_55_43;
	 wire frontend_0_n_55_44;
	 wire frontend_0_n_55_45;
	 wire frontend_0_n_55_46;
	 wire frontend_0_n_55_47;
	 wire frontend_0_n_55_48;
	 wire frontend_0_n_55_49;
	 wire frontend_0_n_55_50;
	 wire frontend_0_n_55_51;
	 wire frontend_0_n_55_52;
	 wire frontend_0_n_55_53;
	 wire frontend_0_n_55_54;
	 wire frontend_0_n_55_55;
	 wire frontend_0_n_55_56;
	 wire frontend_0_n_55_57;
	 wire frontend_0_n_55_58;
	 wire frontend_0_n_55_59;
	 wire frontend_0_n_55_60;
	 wire frontend_0_n_55_61;
	 wire frontend_0_n_55_62;
	 wire frontend_0_n_55_63;
	 wire frontend_0_n_55_64;
	 wire frontend_0_n_55_65;
	 wire frontend_0_n_55_66;
	 wire frontend_0_n_55_67;
	 wire frontend_0_n_55_68;
	 wire frontend_0_n_58_0;
	 wire frontend_0_n_58_1;
	 wire frontend_0_n_58_2;
	 wire frontend_0_n_58_3;
	 wire frontend_0_n_59_0;
	 wire frontend_0_n_59_1;
	 wire frontend_0_n_59_2;
	 wire frontend_0_n_59_3;
	 wire frontend_0_n_59_4;
	 wire frontend_0_n_59_5;
	 wire frontend_0_n_59_6;
	 wire frontend_0_n_60_0;
	 wire frontend_0_irq_detect;
	 wire frontend_0_decode;
	 wire frontend_0_n_64_0;
	 wire [1:0]frontend_0_inst_sz_nxt;
	 wire [1:0]frontend_0_inst_sz;
	 wire frontend_0_n_70_0;
	 wire frontend_0_n_71_0;
	 wire frontend_0_n_72_0;
	 wire frontend_0_n_73_0;
	 wire frontend_0_n_73_1;
	 wire frontend_0_n_73_2;
	 wire frontend_0_n_73_3;
	 wire frontend_0_n_74_0;
	 wire frontend_0_n_75_0;
	 wire frontend_0_n_76_0;
	 wire frontend_0_n_76_1;
	 wire frontend_0_n_76_2;
	 wire frontend_0_n_76_3;
	 wire frontend_0_n_76_4;
	 wire frontend_0_n_76_5;
	 wire frontend_0_n_76_6;
	 wire frontend_0_n_76_7;
	 wire [2:0]frontend_0_i_state_nxt_reg;
	 wire frontend_0_n_76_8;
	 wire frontend_0_n_76_9;
	 wire frontend_0_n_76_10;
	 wire frontend_0_n_76_11;
	 wire frontend_0_n_76_12;
	 wire frontend_0_n_76_13;
	 wire frontend_0_n_76_14;
	 wire frontend_0_n_80_0;
	 wire frontend_0_n_82_0;
	 wire frontend_0_n_82_1;
	 wire frontend_0_n_82_2;
	 wire frontend_0_n_82_3;
	 wire frontend_0_n_82_4;
	 wire frontend_0_n_82_5;
	 wire frontend_0_n_82_6;
	 wire frontend_0_n_82_7;
	 wire frontend_0_n_82_8;
	 wire frontend_0_n_82_9;
	 wire frontend_0_n_82_10;
	 wire [11:0]frontend_0_inst_to_nxt;
	 wire frontend_0_alu_inc;
	 wire [11:0]frontend_0_inst_alu_nxt;
	 wire frontend_0_n_88_0;
	 wire frontend_0_n_88_1;
	 wire frontend_0_n_91_0;
	 wire [3:0]frontend_0_inst_dest_bin;
	 wire frontend_0_n_94_0;
	 wire frontend_0_n_94_1;
	 wire frontend_0_n_94_2;
	 wire frontend_0_n_94_3;
	 wire frontend_0_n_94_4;
	 wire frontend_0_n_94_5;
	 wire frontend_0_n_94_6;
	 wire frontend_0_n_94_7;
	 wire frontend_0_n_94_8;
	 wire frontend_0_n_94_9;
	 wire frontend_0_n_94_10;
	 wire frontend_0_n_94_11;
	 wire frontend_0_n_95_0;
	 wire frontend_0_n_95_1;
	 wire frontend_0_n_95_2;
	 wire frontend_0_n_95_3;
	 wire frontend_0_n_95_4;
	 wire frontend_0_n_95_5;
	 wire frontend_0_n_95_6;
	 wire frontend_0_n_95_7;
	 wire frontend_0_n_95_8;
	 wire frontend_0_n_95_9;
	 wire frontend_0_n_95_10;
	 wire frontend_0_n_95_11;
	 wire frontend_0_n_97_0;
	 wire frontend_0_n_97_1;
	 wire frontend_0_n_97_2;
	 wire frontend_0_n_97_3;
	 wire frontend_0_n_97_4;
	 wire frontend_0_n_97_5;
	 wire frontend_0_n_97_6;
	 wire frontend_0_n_97_7;
	 wire frontend_0_n_97_8;
	 wire frontend_0_n_97_9;
	 wire frontend_0_n_97_10;
	 wire frontend_0_n_97_11;
	 wire frontend_0_n_97_12;
	 wire frontend_0_n_97_13;
	 wire frontend_0_n_97_14;
	 wire frontend_0_n_97_15;
	 wire frontend_0_n_97_16;
	 wire frontend_0_n_97_17;
	 wire frontend_0_n_97_18;
	 wire frontend_0_n_97_19;
	 wire frontend_0_n_98_0;
	 wire frontend_0_n_98_1;
	 wire frontend_0_n_98_2;
	 wire frontend_0_n_98_3;
	 wire frontend_0_n_98_4;
	 wire frontend_0_n_99_0;
	 wire [15:0]frontend_0_ext_nxt;
	 wire frontend_0_n_99_1;
	 wire frontend_0_n_99_2;
	 wire frontend_0_n_99_3;
	 wire frontend_0_n_99_4;
	 wire frontend_0_n_99_5;
	 wire frontend_0_n_99_6;
	 wire frontend_0_n_99_7;
	 wire frontend_0_n_99_8;
	 wire frontend_0_n_99_9;
	 wire frontend_0_n_99_10;
	 wire frontend_0_n_99_11;
	 wire frontend_0_n_99_12;
	 wire frontend_0_n_99_13;
	 wire frontend_0_n_99_14;
	 wire frontend_0_n_99_15;
	 wire frontend_0_n_99_16;
	 wire frontend_0_n_99_17;
	 wire frontend_0_n_101_0;
	 wire frontend_0_n_101_1;
	 wire [2:0]frontend_0_inst_jmp_bin;
	 wire frontend_0_n_105_0;
	 wire frontend_0_n_105_1;
	 wire frontend_0_n_105_2;
	 wire frontend_0_n_105_3;
	 wire frontend_0_n_105_4;
	 wire frontend_0_n_105_5;
	 wire frontend_0_n_105_6;
	 wire frontend_0_n_110_0;
	 wire frontend_0_n_110_1;
	 wire frontend_0_n_110_2;
	 wire frontend_0_n_110_3;
	 wire frontend_0_n_110_4;
	 wire frontend_0_n_110_5;
	 wire frontend_0_n_110_6;
	 wire frontend_0_n_110_7;
	 wire frontend_0_n_110_8;
	 wire frontend_0_n_110_9;
	 wire frontend_0_n_110_10;
	 wire frontend_0_n_110_11;
	 wire frontend_0_n_110_12;
	 wire frontend_0_n_110_13;
	 wire frontend_0_n_110_14;
	 wire frontend_0_n_110_15;
	 wire frontend_0_n_110_16;
	 wire frontend_0_n_110_17;
	 wire frontend_0_n_110_18;
	 wire frontend_0_n_110_19;
	 wire frontend_0_n_110_20;
	 wire frontend_0_n_110_21;
	 wire frontend_0_n_110_22;
	 wire frontend_0_n_110_23;
	 wire frontend_0_n_110_24;
	 wire frontend_0_n_110_25;
	 wire frontend_0_n_110_26;
	 wire frontend_0_n_110_27;
	 wire frontend_0_n_110_28;
	 wire frontend_0_n_110_29;
	 wire frontend_0_n_110_30;
	 wire frontend_0_n_110_31;
	 wire frontend_0_n_110_32;
	 wire frontend_0_n_110_33;
	 wire frontend_0_n_110_34;
	 wire frontend_0_n_110_35;
	 wire frontend_0_n_111_0;
	 wire frontend_0_n_111_1;
	 wire frontend_0_n_111_2;
	 wire frontend_0_n_111_3;
	 wire frontend_0_n_111_4;
	 wire [3:0]frontend_0_inst_src_bin;
	 wire frontend_0_n_114_0;
	 wire frontend_0_n_114_1;
	 wire frontend_0_n_114_2;
	 wire frontend_0_n_114_3;
	 wire frontend_0_n_114_4;
	 wire frontend_0_n_114_5;
	 wire frontend_0_n_114_6;
	 wire frontend_0_n_114_7;
	 wire frontend_0_n_114_8;
	 wire frontend_0_n_114_9;
	 wire frontend_0_n_114_10;
	 wire frontend_0_n_114_11;
	 wire frontend_0_n_115_0;
	 wire frontend_0_n_115_1;
	 wire frontend_0_n_115_2;
	 wire frontend_0_n_115_3;
	 wire frontend_0_n_115_4;
	 wire frontend_0_n_115_5;
	 wire frontend_0_n_115_6;
	 wire frontend_0_n_115_7;
	 wire frontend_0_n_115_8;
	 wire frontend_0_n_115_9;
	 wire frontend_0_n_115_10;
	 wire frontend_0_n_115_11;
	 wire frontend_0_n_115_12;
	 wire frontend_0_n_115_13;
	 wire frontend_0_n_115_14;
	 wire frontend_0_n_115_15;
	 wire frontend_0_n_115_16;
	 wire frontend_0_n_115_17;
	 wire frontend_0_n_115_18;
	 wire frontend_0_n_115_19;
	 wire [5:0]frontend_0_irq_num;
	 wire frontend_0_n_118_0;
	 wire frontend_0_n_118_1;
	 wire frontend_0_n_118_2;
	 wire frontend_0_n_118_3;
	 wire frontend_0_n_118_4;
	 wire frontend_0_n_118_5;
	 wire frontend_0_n_118_6;
	 wire frontend_0_n_118_7;
	 wire frontend_0_n_118_8;
	 wire frontend_0_n_118_9;
	 wire frontend_0_n_118_10;
	 wire frontend_0_n_118_11;
	 wire frontend_0_n_118_12;
	 wire frontend_0_n_118_13;
	 wire frontend_0_n_118_14;
	 wire frontend_0_n_118_15;
	 wire frontend_0_n_118_16;
	 wire frontend_0_n_118_17;
	 wire frontend_0_n_118_18;
	 wire frontend_0_n_118_19;
	 wire frontend_0_n_118_20;
	 wire frontend_0_n_118_21;
	 wire frontend_0_n_118_22;
	 wire frontend_0_n_118_23;
	 wire frontend_0_n_118_24;
	 wire frontend_0_n_118_25;
	 wire frontend_0_n_118_26;
	 wire frontend_0_n_118_27;
	 wire frontend_0_n_118_28;
	 wire frontend_0_n_118_29;
	 wire frontend_0_n_118_30;
	 wire frontend_0_n_118_31;
	 wire frontend_0_n_118_32;
	 wire frontend_0_n_118_33;
	 wire frontend_0_n_118_34;
	 wire frontend_0_n_118_35;
	 wire frontend_0_n_118_36;
	 wire frontend_0_n_118_37;
	 wire frontend_0_n_118_38;
	 wire frontend_0_n_118_39;
	 wire frontend_0_n_118_40;
	 wire frontend_0_n_118_41;
	 wire frontend_0_n_118_42;
	 wire frontend_0_n_118_43;
	 wire frontend_0_n_118_44;
	 wire frontend_0_n_118_45;
	 wire frontend_0_n_118_46;
	 wire frontend_0_n_118_47;
	 wire frontend_0_n_118_48;
	 wire frontend_0_n_118_49;
	 wire frontend_0_n_118_50;
	 wire frontend_0_n_118_51;
	 wire frontend_0_n_118_52;
	 wire frontend_0_n_118_53;
	 wire frontend_0_n_118_54;
	 wire frontend_0_n_118_55;
	 wire frontend_0_n_118_56;
	 wire frontend_0_n_120_0;
	 wire frontend_0_n_120_1;
	 wire frontend_0_n_120_2;
	 wire frontend_0_n_120_3;
	 wire frontend_0_n_120_4;
	 wire frontend_0_n_120_5;
	 wire frontend_0_n_120_6;
	 wire frontend_0_n_120_7;
	 wire frontend_0_n_120_8;
	 wire frontend_0_n_120_9;
	 wire frontend_0_n_120_10;
	 wire frontend_0_n_120_11;
	 wire frontend_0_n_120_12;
	 wire frontend_0_n_120_13;
	 wire frontend_0_n_120_14;
	 wire frontend_0_n_120_15;
	 wire frontend_0_n_120_16;
	 wire frontend_0_n_120_17;
	 wire frontend_0_n_120_18;
	 wire frontend_0_n_120_19;
	 wire frontend_0_n_120_20;
	 wire frontend_0_n_122_0;
	 wire frontend_0_n_122_1;
	 wire frontend_0_n_122_2;
	 wire frontend_0_fetch;
	 wire [15:0]frontend_0_pc_incr;
	 wire frontend_0_n_124_0;
	 wire frontend_0_n_124_1;
	 wire frontend_0_n_124_2;
	 wire frontend_0_n_124_3;
	 wire frontend_0_n_124_4;
	 wire frontend_0_n_124_5;
	 wire frontend_0_n_124_6;
	 wire frontend_0_n_124_7;
	 wire frontend_0_n_124_8;
	 wire frontend_0_n_124_9;
	 wire frontend_0_n_124_10;
	 wire frontend_0_n_124_11;
	 wire frontend_0_n_124_12;
	 wire frontend_0_n_124_13;
	 wire frontend_0_n_124_14;
	 wire frontend_0_n_125_0;
	 wire frontend_0_n_126_0;
	 wire frontend_0_n_126_1;
	 wire frontend_0_n_126_2;
	 wire frontend_0_n_126_3;
	 wire frontend_0_n_126_4;
	 wire frontend_0_n_126_5;
	 wire frontend_0_n_126_6;
	 wire frontend_0_n_126_7;
	 wire frontend_0_n_126_8;
	 wire frontend_0_n_126_9;
	 wire frontend_0_n_126_10;
	 wire frontend_0_n_126_11;
	 wire frontend_0_n_126_12;
	 wire frontend_0_n_126_13;
	 wire frontend_0_n_126_14;
	 wire frontend_0_n_126_15;
	 wire frontend_0_n_127_0;
	 wire frontend_0_n_127_1;
	 wire frontend_0_n_127_2;
	 wire frontend_0_n_127_3;
	 wire frontend_0_n_127_4;
	 wire frontend_0_n_127_5;
	 wire frontend_0_n_127_6;
	 wire frontend_0_n_127_7;
	 wire frontend_0_n_127_8;
	 wire frontend_0_n_127_9;
	 wire frontend_0_n_127_10;
	 wire frontend_0_n_127_11;
	 wire frontend_0_n_127_12;
	 wire frontend_0_n_127_13;
	 wire frontend_0_n_127_14;
	 wire frontend_0_n_127_15;
	 wire frontend_0_n_127_16;
	 wire frontend_0_pmem_busy;
	 wire frontend_0_n_128_0;
	 wire frontend_0_n_128_1;
	 wire frontend_0_n_130_0;
	 wire frontend_0_n_130_1;
	 wire frontend_0_n_130_2;
	 wire frontend_0_n_130_3;
	 wire frontend_0_n_91;
	 wire frontend_0_n_0;
	 wire frontend_0_n_87;
	 wire frontend_0_n_1;
	 wire frontend_0_n_2;
	 wire frontend_0_n_3;
	 wire frontend_0_n_88;
	 wire frontend_0_n_89;
	 wire frontend_0_n_5;
	 wire frontend_0_n_55;
	 wire frontend_0_n_10;
	 wire frontend_0_n_29;
	 wire frontend_0_n_37;
	 wire frontend_0_n_28;
	 wire frontend_0_n_36;
	 wire frontend_0_n_9;
	 wire frontend_0_n_49;
	 wire frontend_0_n_17;
	 wire frontend_0_n_18;
	 wire frontend_0_n_48;
	 wire frontend_0_n_4;
	 wire frontend_0_n_67;
	 wire frontend_0_n_73;
	 wire frontend_0_n_51;
	 wire frontend_0_n_52;
	 wire frontend_0_n_50;
	 wire frontend_0_n_11;
	 wire frontend_0_n_43;
	 wire frontend_0_n_68;
	 wire frontend_0_n_45;
	 wire frontend_0_n_69;
	 wire frontend_0_n_70;
	 wire frontend_0_n_46;
	 wire frontend_0_n_47;
	 wire frontend_0_n_44;
	 wire frontend_0_n_72;
	 wire frontend_0_n_71;
	 wire frontend_0_n_56;
	 wire frontend_0_n_54;
	 wire frontend_0_n_20;
	 wire frontend_0_n_19;
	 wire frontend_0_n_26;
	 wire frontend_0_n_34;
	 wire frontend_0_n_27;
	 wire frontend_0_n_35;
	 wire frontend_0_n_53;
	 wire frontend_0_n_58;
	 wire frontend_0_n_6;
	 wire frontend_0_n_12;
	 wire frontend_0_n_38;
	 wire frontend_0_n_39;
	 wire frontend_0_n_62;
	 wire frontend_0_n_21;
	 wire frontend_0_n_63;
	 wire frontend_0_n_64;
	 wire frontend_0_n_57;
	 wire frontend_0_n_13;
	 wire frontend_0_n_7;
	 wire frontend_0_n_15;
	 wire frontend_0_n_16;
	 wire frontend_0_n_14;
	 wire frontend_0_n_61;
	 wire frontend_0_n_66;
	 wire frontend_0_n_65;
	 wire frontend_0_n_41;
	 wire frontend_0_n_42;
	 wire frontend_0_n_40;
	 wire frontend_0_n_59;
	 wire frontend_0_n_60;
	 wire frontend_0_n_82;
	 wire frontend_0_n_83;
	 wire frontend_0_n_86;
	 wire frontend_0_n_74;
	 wire frontend_0_n_75;
	 wire frontend_0_n_76;
	 wire frontend_0_n_79;
	 wire frontend_0_n_80;
	 wire frontend_0_n_90;
	 wire frontend_0_n_85;
	 wire frontend_0_n_81;
	 wire frontend_0_n_77;
	 wire frontend_0_n_78;
	 wire frontend_0_n_84;
	 wire frontend_0_n_92;
	 wire frontend_0_n_98;
	 wire frontend_0_n_100;
	 wire frontend_0_n_108;
	 wire frontend_0_n_24;
	 wire frontend_0_n_32;
	 wire frontend_0_n_22;
	 wire frontend_0_n_30;
	 wire frontend_0_n_104;
	 wire frontend_0_n_107;
	 wire frontend_0_n_25;
	 wire frontend_0_n_33;
	 wire frontend_0_n_94;
	 wire frontend_0_n_97;
	 wire frontend_0_n_96;
	 wire frontend_0_n_95;
	 wire frontend_0_n_105;
	 wire frontend_0_n_106;
	 wire frontend_0_n_103;
	 wire frontend_0_n_99;
	 wire frontend_0_n_102;
	 wire frontend_0_n_101;
	 wire frontend_0_n_110;
	 wire frontend_0_n_109;
	 wire frontend_0_n_144;
	 wire frontend_0_n_111;
	 wire frontend_0_n_127;
	 wire frontend_0_n_143;
	 wire frontend_0_n_126;
	 wire frontend_0_n_142;
	 wire frontend_0_n_125;
	 wire frontend_0_n_141;
	 wire frontend_0_n_124;
	 wire frontend_0_n_140;
	 wire frontend_0_n_123;
	 wire frontend_0_n_139;
	 wire frontend_0_n_122;
	 wire frontend_0_n_138;
	 wire frontend_0_n_121;
	 wire frontend_0_n_137;
	 wire frontend_0_n_120;
	 wire frontend_0_n_136;
	 wire frontend_0_n_119;
	 wire frontend_0_n_135;
	 wire frontend_0_n_118;
	 wire frontend_0_n_134;
	 wire frontend_0_n_117;
	 wire frontend_0_n_133;
	 wire frontend_0_n_116;
	 wire frontend_0_n_132;
	 wire frontend_0_n_115;
	 wire frontend_0_n_131;
	 wire frontend_0_n_114;
	 wire frontend_0_n_130;
	 wire frontend_0_n_113;
	 wire frontend_0_n_129;
	 wire frontend_0_n_112;
	 wire frontend_0_n_128;
	 wire frontend_0_n_145;
	 wire frontend_0_n_147;
	 wire frontend_0_n_146;
	 wire frontend_0_n_148;
	 wire frontend_0_n_149;
	 wire frontend_0_n_157;
	 wire frontend_0_n_156;
	 wire frontend_0_n_155;
	 wire frontend_0_n_154;
	 wire frontend_0_n_153;
	 wire frontend_0_n_152;
	 wire frontend_0_n_151;
	 wire frontend_0_n_150;
	 wire frontend_0_n_93;
	 wire frontend_0_n_158;
	 wire frontend_0_n_179;
	 wire frontend_0_n_180;
	 wire frontend_0_n_163;
	 wire frontend_0_n_178;
	 wire frontend_0_n_177;
	 wire frontend_0_n_176;
	 wire frontend_0_n_175;
	 wire frontend_0_n_174;
	 wire frontend_0_n_173;
	 wire frontend_0_n_172;
	 wire frontend_0_n_171;
	 wire frontend_0_n_170;
	 wire frontend_0_n_169;
	 wire frontend_0_n_168;
	 wire frontend_0_n_162;
	 wire frontend_0_n_167;
	 wire frontend_0_n_161;
	 wire frontend_0_n_166;
	 wire frontend_0_n_160;
	 wire frontend_0_n_165;
	 wire frontend_0_n_159;
	 wire frontend_0_n_164;
	 wire frontend_0_n_23;
	 wire frontend_0_n_31;
	 wire frontend_0_n_181;
	 wire frontend_0_n_197;
	 wire frontend_0_n_196;
	 wire frontend_0_n_195;
	 wire frontend_0_n_194;
	 wire frontend_0_n_193;
	 wire frontend_0_n_192;
	 wire frontend_0_n_191;
	 wire frontend_0_n_190;
	 wire frontend_0_n_189;
	 wire frontend_0_n_188;
	 wire frontend_0_n_187;
	 wire frontend_0_n_186;
	 wire frontend_0_n_185;
	 wire frontend_0_n_184;
	 wire frontend_0_n_183;
	 wire frontend_0_n_182;
	 wire frontend_0_n_8;
	 wire frontend_0_n_198;
	 wire frontend_0_n_200;
	 wire frontend_0_n_199;
	 wire frontend_0_n_201;
	 wire frontend_0_n_202;
	 wire frontend_0_n_203;
	 wire frontend_0_n_204;
	 wire frontend_0_n_218;
	 wire frontend_0_n_217;
	 wire frontend_0_n_216;
	 wire frontend_0_n_215;
	 wire frontend_0_n_214;
	 wire frontend_0_n_213;
	 wire frontend_0_n_212;
	 wire frontend_0_n_211;
	 wire frontend_0_n_210;
	 wire frontend_0_n_209;
	 wire frontend_0_n_208;
	 wire frontend_0_n_207;
	 wire frontend_0_n_206;
	 wire frontend_0_n_205;
	 wire frontend_0_n_221;
	 wire frontend_0_n_220;
	 wire frontend_0_n_222;
	 wire frontend_0_n_237;
	 wire frontend_0_n_236;
	 wire frontend_0_n_235;
	 wire frontend_0_n_234;
	 wire frontend_0_n_233;
	 wire frontend_0_n_232;
	 wire frontend_0_n_231;
	 wire frontend_0_n_230;
	 wire frontend_0_n_229;
	 wire frontend_0_n_228;
	 wire frontend_0_n_227;
	 wire frontend_0_n_226;
	 wire frontend_0_n_225;
	 wire frontend_0_n_224;
	 wire frontend_0_n_238;
	 wire frontend_0_n_223;
	 wire frontend_0_n_240;
	 wire frontend_0_n_239;
	 wire frontend_0_n_219;
	 wire [3:0]execution_unit_0_alu_stat_wr;
	 wire [3:0]execution_unit_0_alu_stat;
	 wire [15:0]execution_unit_0_alu_out;
	 wire [3:0]execution_unit_0_status;
	 wire [15:0]execution_unit_0_reg_src;
	 wire execution_unit_0_n_0_0;
	 wire execution_unit_0_n_0_1;
	 wire execution_unit_0_n_0_2;
	 wire execution_unit_0_n_0_3;
	 wire execution_unit_0_reg_sr_clr;
	 wire execution_unit_0_n_4_0;
	 wire execution_unit_0_n_4_1;
	 wire execution_unit_0_mb_wr_det;
	 wire execution_unit_0_n_7_0;
	 wire execution_unit_0_n_7_1;
	 wire execution_unit_0_n_7_2;
	 wire execution_unit_0_n_7_3;
	 wire execution_unit_0_n_7_4;
	 wire execution_unit_0_n_8_0;
	 wire execution_unit_0_n_8_1;
	 wire execution_unit_0_n_8_2;
	 wire execution_unit_0_n_8_3;
	 wire execution_unit_0_mab_lsb;
	 wire [15:0]execution_unit_0_mdb_out_nxt;
	 wire execution_unit_0_n_13_0;
	 wire execution_unit_0_n_13_1;
	 wire execution_unit_0_n_13_2;
	 wire execution_unit_0_n_13_3;
	 wire execution_unit_0_n_13_4;
	 wire execution_unit_0_n_13_5;
	 wire execution_unit_0_n_13_6;
	 wire execution_unit_0_n_13_7;
	 wire execution_unit_0_n_13_8;
	 wire execution_unit_0_n_13_9;
	 wire execution_unit_0_n_13_10;
	 wire execution_unit_0_n_13_11;
	 wire execution_unit_0_n_13_12;
	 wire execution_unit_0_n_13_13;
	 wire execution_unit_0_n_13_14;
	 wire execution_unit_0_n_13_15;
	 wire execution_unit_0_n_13_16;
	 wire execution_unit_0_n_13_17;
	 wire execution_unit_0_n_13_18;
	 wire execution_unit_0_n_14_0;
	 wire execution_unit_0_n_14_1;
	 wire execution_unit_0_n_15_0;
	 wire execution_unit_0_n_15_1;
	 wire execution_unit_0_n_15_2;
	 wire execution_unit_0_n_15_3;
	 wire execution_unit_0_n_17_0;
	 wire execution_unit_0_n_17_1;
	 wire execution_unit_0_n_17_2;
	 wire execution_unit_0_n_17_3;
	 wire execution_unit_0_n_17_4;
	 wire execution_unit_0_n_17_5;
	 wire execution_unit_0_n_17_6;
	 wire execution_unit_0_n_17_7;
	 wire execution_unit_0_n_17_8;
	 wire execution_unit_0_n_21_0;
	 wire execution_unit_0_n_21_1;
	 wire execution_unit_0_n_21_2;
	 wire execution_unit_0_n_21_3;
	 wire execution_unit_0_n_21_4;
	 wire execution_unit_0_reg_dest_wr;
	 wire execution_unit_0_n_23_0;
	 wire execution_unit_0_reg_pc_call;
	 wire execution_unit_0_n_30_0;
	 wire execution_unit_0_n_30_1;
	 wire execution_unit_0_n_30_2;
	 wire execution_unit_0_reg_sp_wr;
	 wire execution_unit_0_reg_sr_wr;
	 wire execution_unit_0_n_32_0;
	 wire execution_unit_0_reg_incr;
	 wire execution_unit_0_n_34_0;
	 wire execution_unit_0_n_34_1;
	 wire execution_unit_0_n_34_2;
	 wire execution_unit_0_n_34_3;
	 wire execution_unit_0_n_34_4;
	 wire execution_unit_0_n_34_5;
	 wire execution_unit_0_n_34_6;
	 wire execution_unit_0_n_34_7;
	 wire execution_unit_0_n_34_8;
	 wire execution_unit_0_n_34_9;
	 wire execution_unit_0_n_34_10;
	 wire execution_unit_0_n_34_11;
	 wire execution_unit_0_n_34_12;
	 wire execution_unit_0_n_34_13;
	 wire execution_unit_0_n_34_14;
	 wire execution_unit_0_n_34_15;
	 wire execution_unit_0_n_34_16;
	 wire execution_unit_0_n_34_17;
	 wire execution_unit_0_n_39_0;
	 wire execution_unit_0_n_39_1;
	 wire execution_unit_0_n_39_2;
	 wire execution_unit_0_n_39_3;
	 wire execution_unit_0_n_39_4;
	 wire execution_unit_0_n_39_5;
	 wire execution_unit_0_n_39_6;
	 wire execution_unit_0_n_39_7;
	 wire execution_unit_0_n_39_8;
	 wire execution_unit_0_n_40_0;
	 wire execution_unit_0_n_40_1;
	 wire execution_unit_0_n_40_2;
	 wire execution_unit_0_n_40_3;
	 wire execution_unit_0_n_40_4;
	 wire execution_unit_0_n_40_5;
	 wire execution_unit_0_n_40_6;
	 wire execution_unit_0_n_41_0;
	 wire execution_unit_0_n_41_1;
	 wire execution_unit_0_n_41_2;
	 wire execution_unit_0_n_41_3;
	 wire execution_unit_0_n_41_4;
	 wire execution_unit_0_n_41_5;
	 wire execution_unit_0_n_41_6;
	 wire execution_unit_0_n_41_7;
	 wire execution_unit_0_n_41_8;
	 wire execution_unit_0_n_41_9;
	 wire execution_unit_0_n_41_10;
	 wire execution_unit_0_n_41_11;
	 wire execution_unit_0_n_41_12;
	 wire execution_unit_0_n_41_13;
	 wire execution_unit_0_n_41_14;
	 wire execution_unit_0_n_41_15;
	 wire execution_unit_0_n_41_16;
	 wire execution_unit_0_n_41_17;
	 wire execution_unit_0_n_41_18;
	 wire execution_unit_0_n_41_19;
	 wire execution_unit_0_n_41_20;
	 wire execution_unit_0_n_41_21;
	 wire execution_unit_0_n_41_22;
	 wire execution_unit_0_n_41_23;
	 wire execution_unit_0_n_41_24;
	 wire execution_unit_0_n_41_25;
	 wire execution_unit_0_n_41_26;
	 wire execution_unit_0_n_41_27;
	 wire execution_unit_0_n_41_28;
	 wire execution_unit_0_n_41_29;
	 wire execution_unit_0_n_41_30;
	 wire execution_unit_0_n_41_31;
	 wire execution_unit_0_n_41_32;
	 wire execution_unit_0_n_41_33;
	 wire execution_unit_0_n_41_34;
	 wire execution_unit_0_n_41_35;
	 wire execution_unit_0_n_41_36;
	 wire execution_unit_0_n_41_37;
	 wire execution_unit_0_n_41_38;
	 wire execution_unit_0_n_41_39;
	 wire execution_unit_0_n_41_40;
	 wire execution_unit_0_n_41_41;
	 wire execution_unit_0_n_41_42;
	 wire execution_unit_0_n_41_43;
	 wire execution_unit_0_n_41_44;
	 wire execution_unit_0_n_41_45;
	 wire execution_unit_0_n_41_46;
	 wire execution_unit_0_n_41_47;
	 wire execution_unit_0_n_41_48;
	 wire execution_unit_0_n_41_49;
	 wire execution_unit_0_n_41_50;
	 wire execution_unit_0_n_41_51;
	 wire execution_unit_0_n_41_52;
	 wire execution_unit_0_n_41_53;
	 wire execution_unit_0_n_41_54;
	 wire execution_unit_0_n_41_55;
	 wire execution_unit_0_n_41_56;
	 wire execution_unit_0_n_41_57;
	 wire execution_unit_0_n_41_58;
	 wire execution_unit_0_n_41_59;
	 wire execution_unit_0_n_41_60;
	 wire execution_unit_0_n_41_61;
	 wire execution_unit_0_n_41_62;
	 wire execution_unit_0_n_41_63;
	 wire execution_unit_0_n_41_64;
	 wire execution_unit_0_n_41_65;
	 wire execution_unit_0_n_41_66;
	 wire execution_unit_0_n_41_67;
	 wire execution_unit_0_n_41_68;
	 wire execution_unit_0_n_41_69;
	 wire execution_unit_0_n_41_70;
	 wire execution_unit_0_n_41_71;
	 wire execution_unit_0_n_41_72;
	 wire execution_unit_0_n_41_73;
	 wire execution_unit_0_n_41_74;
	 wire execution_unit_0_n_41_75;
	 wire execution_unit_0_n_41_76;
	 wire execution_unit_0_n_41_77;
	 wire execution_unit_0_n_41_78;
	 wire execution_unit_0_n_41_79;
	 wire execution_unit_0_mdb_in_buf_en;
	 wire [15:0]execution_unit_0_mdb_in_buf;
	 wire execution_unit_0_mdb_in_buf_valid;
	 wire execution_unit_0_n_44_0;
	 wire execution_unit_0_n_44_1;
	 wire execution_unit_0_n_45_0;
	 wire execution_unit_0_n_45_1;
	 wire execution_unit_0_n_45_2;
	 wire execution_unit_0_n_48_0;
	 wire execution_unit_0_n_48_1;
	 wire execution_unit_0_n_48_2;
	 wire execution_unit_0_n_48_3;
	 wire execution_unit_0_n_48_4;
	 wire execution_unit_0_n_48_5;
	 wire execution_unit_0_n_48_6;
	 wire execution_unit_0_n_48_7;
	 wire execution_unit_0_n_48_8;
	 wire execution_unit_0_n_48_9;
	 wire execution_unit_0_n_49_0;
	 wire execution_unit_0_n_49_1;
	 wire execution_unit_0_n_49_2;
	 wire execution_unit_0_n_49_3;
	 wire execution_unit_0_n_49_4;
	 wire execution_unit_0_n_49_5;
	 wire execution_unit_0_n_49_6;
	 wire execution_unit_0_n_49_7;
	 wire execution_unit_0_n_49_8;
	 wire execution_unit_0_n_49_9;
	 wire execution_unit_0_n_50_0;
	 wire execution_unit_0_n_50_1;
	 wire execution_unit_0_n_50_2;
	 wire execution_unit_0_n_50_3;
	 wire execution_unit_0_n_50_4;
	 wire execution_unit_0_n_50_5;
	 wire execution_unit_0_n_50_6;
	 wire execution_unit_0_n_50_7;
	 wire execution_unit_0_n_50_8;
	 wire execution_unit_0_n_50_9;
	 wire execution_unit_0_n_50_10;
	 wire execution_unit_0_n_50_11;
	 wire execution_unit_0_n_50_12;
	 wire execution_unit_0_n_50_13;
	 wire execution_unit_0_n_50_14;
	 wire execution_unit_0_n_50_15;
	 wire execution_unit_0_n_50_16;
	 wire execution_unit_0_n_50_17;
	 wire execution_unit_0_n_50_18;
	 wire execution_unit_0_n_50_19;
	 wire execution_unit_0_n_50_20;
	 wire execution_unit_0_n_50_21;
	 wire execution_unit_0_n_50_22;
	 wire execution_unit_0_n_50_23;
	 wire execution_unit_0_n_50_24;
	 wire execution_unit_0_n_50_25;
	 wire execution_unit_0_n_50_26;
	 wire execution_unit_0_n_50_27;
	 wire execution_unit_0_n_50_28;
	 wire execution_unit_0_n_50_29;
	 wire execution_unit_0_n_50_30;
	 wire execution_unit_0_n_50_31;
	 wire execution_unit_0_n_50_32;
	 wire execution_unit_0_n_50_33;
	 wire execution_unit_0_n_50_34;
	 wire execution_unit_0_n_50_35;
	 wire execution_unit_0_n_50_36;
	 wire execution_unit_0_n_50_37;
	 wire execution_unit_0_n_50_38;
	 wire execution_unit_0_n_50_39;
	 wire execution_unit_0_n_50_40;
	 wire execution_unit_0_n_50_41;
	 wire execution_unit_0_n_50_42;
	 wire execution_unit_0_n_50_43;
	 wire execution_unit_0_n_50_44;
	 wire execution_unit_0_n_50_45;
	 wire execution_unit_0_n_50_46;
	 wire execution_unit_0_n_50_47;
	 wire execution_unit_0_n_50_48;
	 wire execution_unit_0_n_50_49;
	 wire execution_unit_0_n_50_50;
	 wire execution_unit_0_n_50_51;
	 wire execution_unit_0_n_50_52;
	 wire execution_unit_0_n_50_53;
	 wire execution_unit_0_n_50_54;
	 wire execution_unit_0_n_50_55;
	 wire execution_unit_0_n_50_56;
	 wire execution_unit_0_n_50_57;
	 wire execution_unit_0_n_50_58;
	 wire execution_unit_0_n_50_59;
	 wire execution_unit_0_n_50_60;
	 wire execution_unit_0_n_50_61;
	 wire execution_unit_0_n_50_62;
	 wire execution_unit_0_n_50_63;
	 wire execution_unit_0_n_50_64;
	 wire execution_unit_0_n_50_65;
	 wire execution_unit_0_n_50_66;
	 wire execution_unit_0_n_50_67;
	 wire execution_unit_0_n_50_68;
	 wire execution_unit_0_n_50_69;
	 wire execution_unit_0_n_50_70;
	 wire execution_unit_0_n_50_71;
	 wire execution_unit_0_n_50_72;
	 wire execution_unit_0_n_50_73;
	 wire execution_unit_0_n_50_74;
	 wire execution_unit_0_n_50_75;
	 wire execution_unit_0_n_50_76;
	 wire execution_unit_0_n_50_77;
	 wire execution_unit_0_n_50_78;
	 wire execution_unit_0_n_50_79;
	 wire execution_unit_0_n_50_80;
	 wire execution_unit_0_n_50_81;
	 wire execution_unit_0_n_50_82;
	 wire execution_unit_0_n_50_83;
	 wire execution_unit_0_n_50_84;
	 wire execution_unit_0_n_50_85;
	 wire execution_unit_0_n_50_86;
	 wire execution_unit_0_n_50_87;
	 wire execution_unit_0_n_50_88;
	 wire execution_unit_0_n_50_89;
	 wire execution_unit_0_n_50_90;
	 wire execution_unit_0_n_50_91;
	 wire execution_unit_0_n_50_92;
	 wire execution_unit_0_n_50_93;
	 wire execution_unit_0_n_50_94;
	 wire execution_unit_0_n_50_95;
	 wire execution_unit_0_n_0;
	 wire execution_unit_0_n_69;
	 wire execution_unit_0_n_1;
	 wire execution_unit_0_n_2;
	 wire execution_unit_0_n_73;
	 wire execution_unit_0_n_74;
	 wire execution_unit_0_n_3;
	 wire execution_unit_0_n_40;
	 wire execution_unit_0_n_10;
	 wire execution_unit_0_n_67;
	 wire execution_unit_0_n_68;
	 wire execution_unit_0_n_72;
	 wire execution_unit_0_n_75;
	 wire execution_unit_0_n_47;
	 wire execution_unit_0_n_13;
	 wire execution_unit_0_n_11;
	 wire execution_unit_0_n_6;
	 wire execution_unit_0_n_5;
	 wire execution_unit_0_n_12;
	 wire execution_unit_0_n_4;
	 wire execution_unit_0_n_9;
	 wire execution_unit_0_n_16;
	 wire execution_unit_0_n_18;
	 wire execution_unit_0_n_49;
	 wire execution_unit_0_n_48;
	 wire execution_unit_0_n_65;
	 wire execution_unit_0_n_37;
	 wire execution_unit_0_n_38;
	 wire execution_unit_0_n_71;
	 wire execution_unit_0_n_76;
	 wire execution_unit_0_n_41;
	 wire execution_unit_0_n_42;
	 wire execution_unit_0_n_43;
	 wire execution_unit_0_n_8;
	 wire execution_unit_0_n_44;
	 wire execution_unit_0_n_46;
	 wire execution_unit_0_n_66;
	 wire execution_unit_0_n_7;
	 wire execution_unit_0_n_45;
	 wire execution_unit_0_n_70;
	 wire execution_unit_0_n_77;
	 wire execution_unit_0_n_93;
	 wire execution_unit_0_n_64;
	 wire execution_unit_0_n_92;
	 wire execution_unit_0_n_63;
	 wire execution_unit_0_n_91;
	 wire execution_unit_0_n_62;
	 wire execution_unit_0_n_90;
	 wire execution_unit_0_n_61;
	 wire execution_unit_0_n_89;
	 wire execution_unit_0_n_60;
	 wire execution_unit_0_n_88;
	 wire execution_unit_0_n_59;
	 wire execution_unit_0_n_87;
	 wire execution_unit_0_n_58;
	 wire execution_unit_0_n_86;
	 wire execution_unit_0_n_57;
	 wire execution_unit_0_n_85;
	 wire execution_unit_0_n_56;
	 wire execution_unit_0_n_84;
	 wire execution_unit_0_n_55;
	 wire execution_unit_0_n_83;
	 wire execution_unit_0_n_54;
	 wire execution_unit_0_n_82;
	 wire execution_unit_0_n_53;
	 wire execution_unit_0_n_81;
	 wire execution_unit_0_n_52;
	 wire execution_unit_0_n_80;
	 wire execution_unit_0_n_51;
	 wire execution_unit_0_n_79;
	 wire execution_unit_0_n_50;
	 wire execution_unit_0_n_78;
	 wire execution_unit_0_n_102;
	 wire execution_unit_0_n_98;
	 wire execution_unit_0_n_103;
	 wire execution_unit_0_n_96;
	 wire execution_unit_0_n_97;
	 wire execution_unit_0_n_95;
	 wire execution_unit_0_n_101;
	 wire execution_unit_0_n_105;
	 wire execution_unit_0_n_94;
	 wire execution_unit_0_n_106;
	 wire execution_unit_0_n_39;
	 wire execution_unit_0_n_100;
	 wire execution_unit_0_n_107;
	 wire execution_unit_0_n_99;
	 wire execution_unit_0_n_108;
	 wire execution_unit_0_n_104;
	 wire execution_unit_0_n_124;
	 wire execution_unit_0_n_123;
	 wire execution_unit_0_n_122;
	 wire execution_unit_0_n_121;
	 wire execution_unit_0_n_120;
	 wire execution_unit_0_n_119;
	 wire execution_unit_0_n_118;
	 wire execution_unit_0_n_117;
	 wire execution_unit_0_n_116;
	 wire execution_unit_0_n_115;
	 wire execution_unit_0_n_114;
	 wire execution_unit_0_n_113;
	 wire execution_unit_0_n_112;
	 wire execution_unit_0_n_111;
	 wire execution_unit_0_n_110;
	 wire execution_unit_0_n_109;
	 wire execution_unit_0_n_15;
	 wire execution_unit_0_n_14;
	 wire execution_unit_0_n_34;
	 wire execution_unit_0_n_35;
	 wire execution_unit_0_n_36;
	 wire execution_unit_0_n_17;
	 wire execution_unit_0_n_26;
	 wire execution_unit_0_n_33;
	 wire execution_unit_0_n_25;
	 wire execution_unit_0_n_32;
	 wire execution_unit_0_n_24;
	 wire execution_unit_0_n_31;
	 wire execution_unit_0_n_23;
	 wire execution_unit_0_n_30;
	 wire execution_unit_0_n_22;
	 wire execution_unit_0_n_29;
	 wire execution_unit_0_n_21;
	 wire execution_unit_0_n_28;
	 wire execution_unit_0_n_20;
	 wire execution_unit_0_n_27;
	 wire execution_unit_0_n_19;
	 wire execution_unit_0_alu_0_op_bit8_msk;
	 wire execution_unit_0_alu_0_op_src_inv_cmd;
	 wire execution_unit_0_alu_0_n_4_0;
	 wire execution_unit_0_alu_0_n_4_1;
	 wire execution_unit_0_alu_0_n_4_2;
	 wire execution_unit_0_alu_0_n_4_3;
	 wire execution_unit_0_alu_0_n_4_4;
	 wire execution_unit_0_alu_0_n_4_5;
	 wire [3:0]execution_unit_0_alu_0_X;
	 wire execution_unit_0_alu_0_n_4_6;
	 wire execution_unit_0_alu_0_n_4_7;
	 wire execution_unit_0_alu_0_n_4_8;
	 wire execution_unit_0_alu_0_n_5_0;
	 wire execution_unit_0_alu_0_n_5_1;
	 wire execution_unit_0_alu_0_n_5_2;
	 wire execution_unit_0_alu_0_n_5_3;
	 wire execution_unit_0_alu_0_n_5_4;
	 wire execution_unit_0_alu_0_n_5_5;
	 wire execution_unit_0_alu_0_n_6_0;
	 wire execution_unit_0_alu_0_alu_short_thro;
	 wire execution_unit_0_alu_0_n_7_0;
	 wire execution_unit_0_alu_0_n_7_1;
	 wire execution_unit_0_alu_0_n_7_2;
	 wire execution_unit_0_alu_0_n_7_3;
	 wire execution_unit_0_alu_0_n_7_4;
	 wire execution_unit_0_alu_0_n_7_5;
	 wire execution_unit_0_alu_0_n_7_6;
	 wire execution_unit_0_alu_0_n_7_7;
	 wire execution_unit_0_alu_0_n_7_8;
	 wire execution_unit_0_alu_0_n_7_9;
	 wire execution_unit_0_alu_0_n_7_10;
	 wire execution_unit_0_alu_0_n_7_11;
	 wire execution_unit_0_alu_0_n_7_12;
	 wire execution_unit_0_alu_0_n_7_13;
	 wire execution_unit_0_alu_0_n_7_14;
	 wire execution_unit_0_alu_0_n_7_15;
	 wire execution_unit_0_alu_0_n_7_16;
	 wire execution_unit_0_alu_0_n_7_17;
	 wire execution_unit_0_alu_0_n_7_18;
	 wire execution_unit_0_alu_0_n_7_19;
	 wire execution_unit_0_alu_0_n_7_20;
	 wire execution_unit_0_alu_0_n_7_21;
	 wire execution_unit_0_alu_0_n_7_22;
	 wire execution_unit_0_alu_0_n_7_23;
	 wire execution_unit_0_alu_0_n_7_24;
	 wire execution_unit_0_alu_0_n_7_25;
	 wire execution_unit_0_alu_0_n_7_26;
	 wire execution_unit_0_alu_0_n_7_27;
	 wire execution_unit_0_alu_0_n_7_28;
	 wire execution_unit_0_alu_0_n_7_29;
	 wire execution_unit_0_alu_0_n_7_30;
	 wire execution_unit_0_alu_0_n_7_31;
	 wire execution_unit_0_alu_0_n_7_32;
	 wire execution_unit_0_alu_0_n_7_33;
	 wire execution_unit_0_alu_0_n_7_34;
	 wire execution_unit_0_alu_0_n_7_35;
	 wire execution_unit_0_alu_0_n_7_36;
	 wire execution_unit_0_alu_0_n_7_37;
	 wire execution_unit_0_alu_0_n_7_38;
	 wire execution_unit_0_alu_0_n_7_39;
	 wire execution_unit_0_alu_0_n_7_40;
	 wire execution_unit_0_alu_0_n_7_41;
	 wire execution_unit_0_alu_0_n_7_42;
	 wire execution_unit_0_alu_0_n_7_43;
	 wire execution_unit_0_alu_0_n_7_44;
	 wire execution_unit_0_alu_0_n_7_45;
	 wire execution_unit_0_alu_0_n_7_46;
	 wire execution_unit_0_alu_0_n_7_47;
	 wire execution_unit_0_alu_0_n_7_48;
	 wire execution_unit_0_alu_0_n_7_49;
	 wire execution_unit_0_alu_0_n_7_50;
	 wire execution_unit_0_alu_0_n_7_51;
	 wire execution_unit_0_alu_0_n_7_52;
	 wire execution_unit_0_alu_0_n_7_53;
	 wire execution_unit_0_alu_0_n_7_54;
	 wire execution_unit_0_alu_0_n_7_55;
	 wire execution_unit_0_alu_0_n_7_56;
	 wire execution_unit_0_alu_0_n_7_57;
	 wire execution_unit_0_alu_0_n_7_58;
	 wire execution_unit_0_alu_0_n_7_59;
	 wire execution_unit_0_alu_0_n_7_60;
	 wire execution_unit_0_alu_0_n_7_61;
	 wire execution_unit_0_alu_0_n_7_62;
	 wire execution_unit_0_alu_0_n_7_63;
	 wire execution_unit_0_alu_0_n_7_64;
	 wire execution_unit_0_alu_0_n_7_65;
	 wire execution_unit_0_alu_0_n_7_66;
	 wire execution_unit_0_alu_0_n_7_67;
	 wire execution_unit_0_alu_0_n_7_68;
	 wire execution_unit_0_alu_0_n_7_69;
	 wire execution_unit_0_alu_0_n_7_70;
	 wire execution_unit_0_alu_0_n_7_71;
	 wire execution_unit_0_alu_0_n_7_72;
	 wire execution_unit_0_alu_0_n_7_73;
	 wire execution_unit_0_alu_0_n_7_74;
	 wire execution_unit_0_alu_0_n_7_75;
	 wire execution_unit_0_alu_0_n_7_76;
	 wire execution_unit_0_alu_0_n_7_77;
	 wire execution_unit_0_alu_0_n_7_78;
	 wire execution_unit_0_alu_0_n_7_79;
	 wire execution_unit_0_alu_0_n_7_80;
	 wire execution_unit_0_alu_0_n_7_81;
	 wire execution_unit_0_alu_0_n_7_82;
	 wire execution_unit_0_alu_0_n_7_83;
	 wire execution_unit_0_alu_0_n_7_84;
	 wire execution_unit_0_alu_0_n_7_85;
	 wire execution_unit_0_alu_0_n_7_86;
	 wire execution_unit_0_alu_0_n_7_87;
	 wire execution_unit_0_alu_0_n_7_88;
	 wire execution_unit_0_alu_0_n_7_89;
	 wire execution_unit_0_alu_0_n_7_90;
	 wire execution_unit_0_alu_0_n_7_91;
	 wire execution_unit_0_alu_0_n_7_92;
	 wire execution_unit_0_alu_0_n_7_93;
	 wire execution_unit_0_alu_0_n_7_94;
	 wire execution_unit_0_alu_0_n_7_95;
	 wire execution_unit_0_alu_0_n_7_96;
	 wire execution_unit_0_alu_0_n_7_97;
	 wire execution_unit_0_alu_0_n_7_98;
	 wire execution_unit_0_alu_0_n_7_99;
	 wire execution_unit_0_alu_0_n_7_100;
	 wire execution_unit_0_alu_0_n_7_101;
	 wire execution_unit_0_alu_0_n_7_102;
	 wire execution_unit_0_alu_0_n_7_103;
	 wire execution_unit_0_alu_0_n_7_104;
	 wire execution_unit_0_alu_0_n_7_105;
	 wire execution_unit_0_alu_0_n_7_106;
	 wire execution_unit_0_alu_0_n_7_107;
	 wire execution_unit_0_alu_0_n_7_108;
	 wire execution_unit_0_alu_0_n_7_109;
	 wire execution_unit_0_alu_0_n_7_110;
	 wire execution_unit_0_alu_0_n_7_111;
	 wire execution_unit_0_alu_0_n_7_112;
	 wire execution_unit_0_alu_0_n_7_113;
	 wire execution_unit_0_alu_0_n_7_114;
	 wire execution_unit_0_alu_0_n_7_115;
	 wire execution_unit_0_alu_0_n_7_116;
	 wire execution_unit_0_alu_0_n_7_117;
	 wire execution_unit_0_alu_0_n_7_118;
	 wire execution_unit_0_alu_0_n_7_119;
	 wire execution_unit_0_alu_0_n_7_120;
	 wire execution_unit_0_alu_0_n_7_121;
	 wire execution_unit_0_alu_0_n_7_122;
	 wire execution_unit_0_alu_0_n_7_123;
	 wire execution_unit_0_alu_0_n_7_124;
	 wire execution_unit_0_alu_0_n_7_125;
	 wire execution_unit_0_alu_0_n_7_126;
	 wire execution_unit_0_alu_0_n_7_127;
	 wire execution_unit_0_alu_0_n_7_128;
	 wire execution_unit_0_alu_0_n_7_129;
	 wire execution_unit_0_alu_0_n_7_130;
	 wire execution_unit_0_alu_0_n_7_131;
	 wire execution_unit_0_alu_0_n_7_132;
	 wire execution_unit_0_alu_0_n_7_133;
	 wire execution_unit_0_alu_0_n_7_134;
	 wire execution_unit_0_alu_0_n_7_135;
	 wire execution_unit_0_alu_0_n_8_0;
	 wire execution_unit_0_alu_0_n_9_0;
	 wire execution_unit_0_alu_0_n_9_1;
	 wire execution_unit_0_alu_0_n_9_2;
	 wire execution_unit_0_alu_0_n_9_3;
	 wire execution_unit_0_alu_0_n_9_4;
	 wire execution_unit_0_alu_0_n_9_5;
	 wire execution_unit_0_alu_0_n_9_6;
	 wire execution_unit_0_alu_0_n_9_7;
	 wire execution_unit_0_alu_0_n_9_8;
	 wire execution_unit_0_alu_0_n_9_9;
	 wire execution_unit_0_alu_0_n_11_0;
	 wire execution_unit_0_alu_0_n_11_1;
	 wire execution_unit_0_alu_0_n_11_2;
	 wire execution_unit_0_alu_0_n_12_0;
	 wire [4:0]execution_unit_0_alu_0_bcd_add;
	 wire execution_unit_0_alu_0_n_12_1;
	 wire execution_unit_0_alu_0_n_12_2;
	 wire execution_unit_0_alu_0_n_12_3;
	 wire execution_unit_0_alu_0_n_12_4;
	 wire execution_unit_0_alu_0_n_12_5;
	 wire execution_unit_0_alu_0_n_12_6;
	 wire execution_unit_0_alu_0_n_12_7;
	 wire execution_unit_0_alu_0_n_12_8;
	 wire execution_unit_0_alu_0_n_13_0;
	 wire execution_unit_0_alu_0_n_14_0;
	 wire execution_unit_0_alu_0_n_14_1;
	 wire execution_unit_0_alu_0_n_14_2;
	 wire execution_unit_0_alu_0_n_14_3;
	 wire execution_unit_0_alu_0_n_14_4;
	 wire execution_unit_0_alu_0_n_14_5;
	 wire execution_unit_0_alu_0_n_14_6;
	 wire execution_unit_0_alu_0_n_14_7;
	 wire execution_unit_0_alu_0_n_14_8;
	 wire execution_unit_0_alu_0_n_14_9;
	 wire execution_unit_0_alu_0_n_16_0;
	 wire execution_unit_0_alu_0_n_16_1;
	 wire execution_unit_0_alu_0_n_16_2;
	 wire execution_unit_0_alu_0_n_17_0;
	 wire [4:0]execution_unit_0_alu_0_bcd_add0;
	 wire execution_unit_0_alu_0_n_17_1;
	 wire execution_unit_0_alu_0_n_17_2;
	 wire execution_unit_0_alu_0_n_17_3;
	 wire execution_unit_0_alu_0_n_17_4;
	 wire execution_unit_0_alu_0_n_17_5;
	 wire execution_unit_0_alu_0_n_17_6;
	 wire execution_unit_0_alu_0_n_17_7;
	 wire execution_unit_0_alu_0_n_17_8;
	 wire execution_unit_0_alu_0_n_18_0;
	 wire execution_unit_0_alu_0_n_19_0;
	 wire execution_unit_0_alu_0_n_19_1;
	 wire execution_unit_0_alu_0_n_19_2;
	 wire execution_unit_0_alu_0_n_19_3;
	 wire execution_unit_0_alu_0_n_19_4;
	 wire execution_unit_0_alu_0_n_19_5;
	 wire execution_unit_0_alu_0_n_19_6;
	 wire execution_unit_0_alu_0_n_19_7;
	 wire execution_unit_0_alu_0_n_19_8;
	 wire execution_unit_0_alu_0_n_19_9;
	 wire execution_unit_0_alu_0_n_21_0;
	 wire execution_unit_0_alu_0_n_21_1;
	 wire execution_unit_0_alu_0_n_21_2;
	 wire execution_unit_0_alu_0_n_22_0;
	 wire [4:0]execution_unit_0_alu_0_bcd_add1;
	 wire execution_unit_0_alu_0_n_22_1;
	 wire execution_unit_0_alu_0_n_22_2;
	 wire execution_unit_0_alu_0_n_22_3;
	 wire execution_unit_0_alu_0_n_22_4;
	 wire execution_unit_0_alu_0_n_22_5;
	 wire execution_unit_0_alu_0_n_22_6;
	 wire execution_unit_0_alu_0_n_22_7;
	 wire execution_unit_0_alu_0_n_22_8;
	 wire execution_unit_0_alu_0_n_23_0;
	 wire execution_unit_0_alu_0_n_24_0;
	 wire execution_unit_0_alu_0_n_24_1;
	 wire execution_unit_0_alu_0_n_24_2;
	 wire execution_unit_0_alu_0_n_24_3;
	 wire execution_unit_0_alu_0_n_24_4;
	 wire execution_unit_0_alu_0_n_24_5;
	 wire execution_unit_0_alu_0_n_24_6;
	 wire execution_unit_0_alu_0_n_24_7;
	 wire execution_unit_0_alu_0_n_24_8;
	 wire execution_unit_0_alu_0_n_24_9;
	 wire execution_unit_0_alu_0_n_26_0;
	 wire execution_unit_0_alu_0_n_26_1;
	 wire execution_unit_0_alu_0_n_26_2;
	 wire execution_unit_0_alu_0_n_27_0;
	 wire [4:0]execution_unit_0_alu_0_bcd_add2;
	 wire execution_unit_0_alu_0_n_27_1;
	 wire execution_unit_0_alu_0_n_27_2;
	 wire execution_unit_0_alu_0_n_27_3;
	 wire execution_unit_0_alu_0_n_27_4;
	 wire execution_unit_0_alu_0_n_27_5;
	 wire execution_unit_0_alu_0_n_27_6;
	 wire execution_unit_0_alu_0_n_27_7;
	 wire execution_unit_0_alu_0_n_27_8;
	 wire execution_unit_0_alu_0_n_28_0;
	 wire execution_unit_0_alu_0_n_28_1;
	 wire execution_unit_0_alu_0_alu_inc;
	 wire execution_unit_0_alu_0_n_30_0;
	 wire execution_unit_0_alu_0_n_30_1;
	 wire execution_unit_0_alu_0_n_30_2;
	 wire execution_unit_0_alu_0_n_30_3;
	 wire execution_unit_0_alu_0_n_30_4;
	 wire execution_unit_0_alu_0_n_30_5;
	 wire execution_unit_0_alu_0_n_30_6;
	 wire execution_unit_0_alu_0_n_30_7;
	 wire execution_unit_0_alu_0_n_30_8;
	 wire execution_unit_0_alu_0_n_30_9;
	 wire execution_unit_0_alu_0_n_40_0;
	 wire execution_unit_0_alu_0_n_40_1;
	 wire execution_unit_0_alu_0_n_40_2;
	 wire execution_unit_0_alu_0_n_40_3;
	 wire execution_unit_0_alu_0_n_40_4;
	 wire execution_unit_0_alu_0_n_40_5;
	 wire execution_unit_0_alu_0_n_40_6;
	 wire execution_unit_0_alu_0_n_40_7;
	 wire execution_unit_0_alu_0_n_40_8;
	 wire execution_unit_0_alu_0_n_40_9;
	 wire execution_unit_0_alu_0_n_40_10;
	 wire execution_unit_0_alu_0_n_40_11;
	 wire execution_unit_0_alu_0_n_40_12;
	 wire execution_unit_0_alu_0_n_40_13;
	 wire execution_unit_0_alu_0_n_40_14;
	 wire [16:0]execution_unit_0_alu_0_alu_add;
	 wire [16:0]execution_unit_0_alu_0_alu_add_inc;
	 wire execution_unit_0_alu_0_n_41_0;
	 wire execution_unit_0_alu_0_n_41_1;
	 wire execution_unit_0_alu_0_n_41_2;
	 wire execution_unit_0_alu_0_n_41_3;
	 wire execution_unit_0_alu_0_n_41_4;
	 wire execution_unit_0_alu_0_n_41_5;
	 wire execution_unit_0_alu_0_n_41_6;
	 wire execution_unit_0_alu_0_n_41_7;
	 wire execution_unit_0_alu_0_n_41_8;
	 wire execution_unit_0_alu_0_n_41_9;
	 wire execution_unit_0_alu_0_n_41_10;
	 wire execution_unit_0_alu_0_n_41_11;
	 wire execution_unit_0_alu_0_n_41_12;
	 wire execution_unit_0_alu_0_n_41_13;
	 wire execution_unit_0_alu_0_n_41_14;
	 wire execution_unit_0_alu_0_n_41_15;
	 wire execution_unit_0_alu_0_n_41_16;
	 wire execution_unit_0_alu_0_n_43_0;
	 wire execution_unit_0_alu_0_n_44_0;
	 wire execution_unit_0_alu_0_n_44_1;
	 wire execution_unit_0_alu_0_n_44_2;
	 wire execution_unit_0_alu_0_n_44_3;
	 wire execution_unit_0_alu_0_n_44_4;
	 wire execution_unit_0_alu_0_n_44_5;
	 wire execution_unit_0_alu_0_n_44_6;
	 wire execution_unit_0_alu_0_n_44_7;
	 wire execution_unit_0_alu_0_n_44_8;
	 wire execution_unit_0_alu_0_n_44_9;
	 wire execution_unit_0_alu_0_n_44_10;
	 wire execution_unit_0_alu_0_n_44_11;
	 wire execution_unit_0_alu_0_n_44_12;
	 wire execution_unit_0_alu_0_n_44_13;
	 wire execution_unit_0_alu_0_n_44_14;
	 wire execution_unit_0_alu_0_n_44_15;
	 wire execution_unit_0_alu_0_n_44_16;
	 wire execution_unit_0_alu_0_n_46_0;
	 wire execution_unit_0_alu_0_n_46_1;
	 wire execution_unit_0_alu_0_n_46_2;
	 wire execution_unit_0_alu_0_n_48_0;
	 wire execution_unit_0_alu_0_n_48_1;
	 wire execution_unit_0_alu_0_n_48_2;
	 wire execution_unit_0_alu_0_n_49_0;
	 wire execution_unit_0_alu_0_n_49_1;
	 wire execution_unit_0_alu_0_n_49_2;
	 wire execution_unit_0_alu_0_n_49_3;
	 wire execution_unit_0_alu_0_n_49_4;
	 wire execution_unit_0_alu_0_n_49_5;
	 wire execution_unit_0_alu_0_n_49_6;
	 wire execution_unit_0_alu_0_n_49_7;
	 wire execution_unit_0_alu_0_n_49_8;
	 wire execution_unit_0_alu_0_n_49_9;
	 wire execution_unit_0_alu_0_Z;
	 wire execution_unit_0_alu_0_n_51_0;
	 wire execution_unit_0_alu_0_n_51_1;
	 wire execution_unit_0_alu_0_n_51_2;
	 wire execution_unit_0_alu_0_n_51_3;
	 wire execution_unit_0_alu_0_n_51_4;
	 wire execution_unit_0_alu_0_n_51_5;
	 wire execution_unit_0_alu_0_n_51_6;
	 wire execution_unit_0_alu_0_n_51_7;
	 wire execution_unit_0_alu_0_n_51_8;
	 wire execution_unit_0_alu_0_n_51_9;
	 wire execution_unit_0_alu_0_n_51_10;
	 wire execution_unit_0_alu_0_n_51_11;
	 wire execution_unit_0_alu_0_n_51_12;
	 wire execution_unit_0_alu_0_n_51_13;
	 wire execution_unit_0_alu_0_n_51_14;
	 wire execution_unit_0_alu_0_n_51_15;
	 wire execution_unit_0_alu_0_n_51_16;
	 wire execution_unit_0_alu_0_n_51_17;
	 wire execution_unit_0_alu_0_n_51_18;
	 wire execution_unit_0_alu_0_n_51_19;
	 wire execution_unit_0_alu_0_n_51_20;
	 wire execution_unit_0_alu_0_n_51_21;
	 wire execution_unit_0_alu_0_n_51_22;
	 wire execution_unit_0_alu_0_n_104;
	 wire execution_unit_0_alu_0_n_7;
	 wire execution_unit_0_alu_0_n_86;
	 wire execution_unit_0_alu_0_n_87;
	 wire execution_unit_0_alu_0_n_103;
	 wire execution_unit_0_alu_0_n_6;
	 wire execution_unit_0_alu_0_n_102;
	 wire execution_unit_0_alu_0_n_5;
	 wire execution_unit_0_alu_0_n_101;
	 wire execution_unit_0_alu_0_n_4;
	 wire execution_unit_0_alu_0_n_100;
	 wire execution_unit_0_alu_0_n_3;
	 wire execution_unit_0_alu_0_n_19;
	 wire execution_unit_0_alu_0_n_99;
	 wire execution_unit_0_alu_0_n_2;
	 wire execution_unit_0_alu_0_n_18;
	 wire execution_unit_0_alu_0_n_98;
	 wire execution_unit_0_alu_0_n_1;
	 wire execution_unit_0_alu_0_n_17;
	 wire execution_unit_0_alu_0_n_97;
	 wire execution_unit_0_alu_0_n_0;
	 wire execution_unit_0_alu_0_n_16;
	 wire execution_unit_0_alu_0_n_96;
	 wire execution_unit_0_alu_0_n_15;
	 wire execution_unit_0_alu_0_n_95;
	 wire execution_unit_0_alu_0_n_14;
	 wire execution_unit_0_alu_0_n_94;
	 wire execution_unit_0_alu_0_n_13;
	 wire execution_unit_0_alu_0_n_93;
	 wire execution_unit_0_alu_0_n_12;
	 wire execution_unit_0_alu_0_n_92;
	 wire execution_unit_0_alu_0_n_11;
	 wire execution_unit_0_alu_0_n_91;
	 wire execution_unit_0_alu_0_n_10;
	 wire execution_unit_0_alu_0_n_90;
	 wire execution_unit_0_alu_0_n_9;
	 wire execution_unit_0_alu_0_n_89;
	 wire execution_unit_0_alu_0_n_8;
	 wire execution_unit_0_alu_0_n_88;
	 wire execution_unit_0_alu_0_n_106;
	 wire execution_unit_0_alu_0_n_68;
	 wire execution_unit_0_alu_0_n_67;
	 wire execution_unit_0_alu_0_n_66;
	 wire execution_unit_0_alu_0_n_65;
	 wire execution_unit_0_alu_0_n_56;
	 wire execution_unit_0_alu_0_n_55;
	 wire execution_unit_0_alu_0_n_54;
	 wire execution_unit_0_alu_0_n_53;
	 wire execution_unit_0_alu_0_n_44;
	 wire execution_unit_0_alu_0_n_43;
	 wire execution_unit_0_alu_0_n_42;
	 wire execution_unit_0_alu_0_n_41;
	 wire execution_unit_0_alu_0_n_38;
	 wire execution_unit_0_alu_0_n_40;
	 wire execution_unit_0_alu_0_n_39;
	 wire execution_unit_0_alu_0_n_45;
	 wire execution_unit_0_alu_0_n_46;
	 wire execution_unit_0_alu_0_n_47;
	 wire execution_unit_0_alu_0_n_48;
	 wire execution_unit_0_alu_0_n_49;
	 wire execution_unit_0_alu_0_n_50;
	 wire execution_unit_0_alu_0_n_52;
	 wire execution_unit_0_alu_0_n_51;
	 wire execution_unit_0_alu_0_n_57;
	 wire execution_unit_0_alu_0_n_58;
	 wire execution_unit_0_alu_0_n_59;
	 wire execution_unit_0_alu_0_n_60;
	 wire execution_unit_0_alu_0_n_61;
	 wire execution_unit_0_alu_0_n_62;
	 wire execution_unit_0_alu_0_n_64;
	 wire execution_unit_0_alu_0_n_63;
	 wire execution_unit_0_alu_0_n_69;
	 wire execution_unit_0_alu_0_n_70;
	 wire execution_unit_0_alu_0_n_71;
	 wire execution_unit_0_alu_0_n_72;
	 wire execution_unit_0_alu_0_n_73;
	 wire execution_unit_0_alu_0_n_74;
	 wire execution_unit_0_alu_0_n_76;
	 wire execution_unit_0_alu_0_n_75;
	 wire execution_unit_0_alu_0_n_78;
	 wire execution_unit_0_alu_0_n_77;
	 wire execution_unit_0_alu_0_n_83;
	 wire execution_unit_0_alu_0_n_80;
	 wire execution_unit_0_alu_0_n_79;
	 wire execution_unit_0_alu_0_n_81;
	 wire execution_unit_0_alu_0_n_82;
	 wire execution_unit_0_alu_0_n_84;
	 wire execution_unit_0_alu_0_n_105;
	 wire execution_unit_0_alu_0_n_20;
	 wire execution_unit_0_alu_0_n_37;
	 wire execution_unit_0_alu_0_n_36;
	 wire execution_unit_0_alu_0_n_35;
	 wire execution_unit_0_alu_0_n_34;
	 wire execution_unit_0_alu_0_n_33;
	 wire execution_unit_0_alu_0_n_32;
	 wire execution_unit_0_alu_0_n_31;
	 wire execution_unit_0_alu_0_n_30;
	 wire execution_unit_0_alu_0_n_21;
	 wire execution_unit_0_alu_0_n_29;
	 wire execution_unit_0_alu_0_n_28;
	 wire execution_unit_0_alu_0_n_27;
	 wire execution_unit_0_alu_0_n_26;
	 wire execution_unit_0_alu_0_n_25;
	 wire execution_unit_0_alu_0_n_24;
	 wire execution_unit_0_alu_0_n_23;
	 wire execution_unit_0_alu_0_n_22;
	 wire execution_unit_0_alu_0_n_108;
	 wire execution_unit_0_alu_0_n_110;
	 wire execution_unit_0_alu_0_n_109;
	 wire execution_unit_0_alu_0_n_111;
	 wire execution_unit_0_alu_0_n_112;
	 wire execution_unit_0_alu_0_n_85;
	 wire execution_unit_0_alu_0_n_107;
	 wire execution_unit_0_register_file_0_n_0_0;
	 wire execution_unit_0_register_file_0_n_1_0;
	 wire execution_unit_0_register_file_0_r2_wr;
	 wire execution_unit_0_register_file_0_n_2_0;
	 wire execution_unit_0_register_file_0_n_2_1;
	 wire [4:0]execution_unit_0_register_file_0_r2_nxt;
	 wire execution_unit_0_register_file_0_n_2_2;
	 wire execution_unit_0_register_file_0_n_2_3;
	 wire execution_unit_0_register_file_0_n_2_4;
	 wire execution_unit_0_register_file_0_n_5_0;
	 wire execution_unit_0_register_file_0_n_5_1;
	 wire execution_unit_0_register_file_0_n_5_2;
	 wire execution_unit_0_register_file_0_n_5_3;
	 wire execution_unit_0_register_file_0_n_5_4;
	 wire execution_unit_0_register_file_0_n_5_5;
	 wire execution_unit_0_register_file_0_n_5_6;
	 wire execution_unit_0_register_file_0_n_5_7;
	 wire execution_unit_0_register_file_0_n_5_8;
	 wire execution_unit_0_register_file_0_n_5_9;
	 wire execution_unit_0_register_file_0_n_5_10;
	 wire execution_unit_0_register_file_0_n_5_11;
	 wire execution_unit_0_register_file_0_n_5_12;
	 wire execution_unit_0_register_file_0_n_5_13;
	 wire execution_unit_0_register_file_0_n_5_14;
	 wire execution_unit_0_register_file_0_n_5_15;
	 wire execution_unit_0_register_file_0_n_5_16;
	 wire execution_unit_0_register_file_0_n_6_0;
	 wire execution_unit_0_register_file_0_n_8_0;
	 wire execution_unit_0_register_file_0_n_9_0;
	 wire execution_unit_0_register_file_0_n_10_0;
	 wire execution_unit_0_register_file_0_inst_src_in;
	 wire execution_unit_0_register_file_0_r1_inc;
	 wire execution_unit_0_register_file_0_r1_wr;
	 wire execution_unit_0_register_file_0_n_13_0;
	 wire execution_unit_0_register_file_0_n_13_1;
	 wire execution_unit_0_register_file_0_n_14_0;
	 wire execution_unit_0_register_file_0_r3_wr;
	 wire [15:0]execution_unit_0_register_file_0_r3;
	 wire execution_unit_0_register_file_0_n_17_0;
	 wire execution_unit_0_register_file_0_r4_inc;
	 wire execution_unit_0_register_file_0_r4_wr;
	 wire execution_unit_0_register_file_0_n_20_0;
	 wire [15:0]execution_unit_0_register_file_0_reg_incr_val;
	 wire execution_unit_0_register_file_0_n_22_0;
	 wire execution_unit_0_register_file_0_n_22_1;
	 wire execution_unit_0_register_file_0_n_22_2;
	 wire execution_unit_0_register_file_0_n_22_3;
	 wire execution_unit_0_register_file_0_n_22_4;
	 wire execution_unit_0_register_file_0_n_22_5;
	 wire execution_unit_0_register_file_0_n_22_6;
	 wire execution_unit_0_register_file_0_n_22_7;
	 wire execution_unit_0_register_file_0_n_22_8;
	 wire execution_unit_0_register_file_0_n_22_9;
	 wire execution_unit_0_register_file_0_n_22_10;
	 wire execution_unit_0_register_file_0_n_22_11;
	 wire execution_unit_0_register_file_0_n_22_12;
	 wire execution_unit_0_register_file_0_n_22_13;
	 wire execution_unit_0_register_file_0_n_22_14;
	 wire execution_unit_0_register_file_0_n_22_15;
	 wire [15:0]execution_unit_0_register_file_0_r4;
	 wire execution_unit_0_register_file_0_n_24_0;
	 wire execution_unit_0_register_file_0_n_24_1;
	 wire execution_unit_0_register_file_0_n_24_2;
	 wire execution_unit_0_register_file_0_n_24_3;
	 wire execution_unit_0_register_file_0_n_24_4;
	 wire execution_unit_0_register_file_0_n_24_5;
	 wire execution_unit_0_register_file_0_n_24_6;
	 wire execution_unit_0_register_file_0_n_24_7;
	 wire execution_unit_0_register_file_0_n_24_8;
	 wire execution_unit_0_register_file_0_n_24_9;
	 wire execution_unit_0_register_file_0_n_24_10;
	 wire execution_unit_0_register_file_0_n_24_11;
	 wire execution_unit_0_register_file_0_n_24_12;
	 wire execution_unit_0_register_file_0_n_24_13;
	 wire execution_unit_0_register_file_0_n_24_14;
	 wire execution_unit_0_register_file_0_n_24_15;
	 wire execution_unit_0_register_file_0_n_24_16;
	 wire execution_unit_0_register_file_0_n_25_0;
	 wire execution_unit_0_register_file_0_n_25_1;
	 wire execution_unit_0_register_file_0_n_27_0;
	 wire execution_unit_0_register_file_0_r5_inc;
	 wire execution_unit_0_register_file_0_r5_wr;
	 wire [15:0]execution_unit_0_register_file_0_r5;
	 wire execution_unit_0_register_file_0_n_31_0;
	 wire execution_unit_0_register_file_0_n_31_1;
	 wire execution_unit_0_register_file_0_n_31_2;
	 wire execution_unit_0_register_file_0_n_31_3;
	 wire execution_unit_0_register_file_0_n_31_4;
	 wire execution_unit_0_register_file_0_n_31_5;
	 wire execution_unit_0_register_file_0_n_31_6;
	 wire execution_unit_0_register_file_0_n_31_7;
	 wire execution_unit_0_register_file_0_n_31_8;
	 wire execution_unit_0_register_file_0_n_31_9;
	 wire execution_unit_0_register_file_0_n_31_10;
	 wire execution_unit_0_register_file_0_n_31_11;
	 wire execution_unit_0_register_file_0_n_31_12;
	 wire execution_unit_0_register_file_0_n_31_13;
	 wire execution_unit_0_register_file_0_n_31_14;
	 wire execution_unit_0_register_file_0_n_31_15;
	 wire execution_unit_0_register_file_0_n_31_16;
	 wire execution_unit_0_register_file_0_n_32_0;
	 wire execution_unit_0_register_file_0_n_32_1;
	 wire execution_unit_0_register_file_0_n_34_0;
	 wire execution_unit_0_register_file_0_r6_inc;
	 wire execution_unit_0_register_file_0_r6_wr;
	 wire [15:0]execution_unit_0_register_file_0_r6;
	 wire execution_unit_0_register_file_0_n_38_0;
	 wire execution_unit_0_register_file_0_n_38_1;
	 wire execution_unit_0_register_file_0_n_38_2;
	 wire execution_unit_0_register_file_0_n_38_3;
	 wire execution_unit_0_register_file_0_n_38_4;
	 wire execution_unit_0_register_file_0_n_38_5;
	 wire execution_unit_0_register_file_0_n_38_6;
	 wire execution_unit_0_register_file_0_n_38_7;
	 wire execution_unit_0_register_file_0_n_38_8;
	 wire execution_unit_0_register_file_0_n_38_9;
	 wire execution_unit_0_register_file_0_n_38_10;
	 wire execution_unit_0_register_file_0_n_38_11;
	 wire execution_unit_0_register_file_0_n_38_12;
	 wire execution_unit_0_register_file_0_n_38_13;
	 wire execution_unit_0_register_file_0_n_38_14;
	 wire execution_unit_0_register_file_0_n_38_15;
	 wire execution_unit_0_register_file_0_n_38_16;
	 wire execution_unit_0_register_file_0_n_39_0;
	 wire execution_unit_0_register_file_0_n_39_1;
	 wire execution_unit_0_register_file_0_n_41_0;
	 wire execution_unit_0_register_file_0_r7_inc;
	 wire execution_unit_0_register_file_0_r7_wr;
	 wire [15:0]execution_unit_0_register_file_0_r7;
	 wire execution_unit_0_register_file_0_n_45_0;
	 wire execution_unit_0_register_file_0_n_45_1;
	 wire execution_unit_0_register_file_0_n_45_2;
	 wire execution_unit_0_register_file_0_n_45_3;
	 wire execution_unit_0_register_file_0_n_45_4;
	 wire execution_unit_0_register_file_0_n_45_5;
	 wire execution_unit_0_register_file_0_n_45_6;
	 wire execution_unit_0_register_file_0_n_45_7;
	 wire execution_unit_0_register_file_0_n_45_8;
	 wire execution_unit_0_register_file_0_n_45_9;
	 wire execution_unit_0_register_file_0_n_45_10;
	 wire execution_unit_0_register_file_0_n_45_11;
	 wire execution_unit_0_register_file_0_n_45_12;
	 wire execution_unit_0_register_file_0_n_45_13;
	 wire execution_unit_0_register_file_0_n_45_14;
	 wire execution_unit_0_register_file_0_n_45_15;
	 wire execution_unit_0_register_file_0_n_45_16;
	 wire execution_unit_0_register_file_0_n_46_0;
	 wire execution_unit_0_register_file_0_n_46_1;
	 wire execution_unit_0_register_file_0_n_48_0;
	 wire execution_unit_0_register_file_0_r8_inc;
	 wire execution_unit_0_register_file_0_r8_wr;
	 wire [15:0]execution_unit_0_register_file_0_r8;
	 wire execution_unit_0_register_file_0_n_52_0;
	 wire execution_unit_0_register_file_0_n_52_1;
	 wire execution_unit_0_register_file_0_n_52_2;
	 wire execution_unit_0_register_file_0_n_52_3;
	 wire execution_unit_0_register_file_0_n_52_4;
	 wire execution_unit_0_register_file_0_n_52_5;
	 wire execution_unit_0_register_file_0_n_52_6;
	 wire execution_unit_0_register_file_0_n_52_7;
	 wire execution_unit_0_register_file_0_n_52_8;
	 wire execution_unit_0_register_file_0_n_52_9;
	 wire execution_unit_0_register_file_0_n_52_10;
	 wire execution_unit_0_register_file_0_n_52_11;
	 wire execution_unit_0_register_file_0_n_52_12;
	 wire execution_unit_0_register_file_0_n_52_13;
	 wire execution_unit_0_register_file_0_n_52_14;
	 wire execution_unit_0_register_file_0_n_52_15;
	 wire execution_unit_0_register_file_0_n_52_16;
	 wire execution_unit_0_register_file_0_n_53_0;
	 wire execution_unit_0_register_file_0_n_53_1;
	 wire execution_unit_0_register_file_0_n_55_0;
	 wire execution_unit_0_register_file_0_r9_inc;
	 wire execution_unit_0_register_file_0_r9_wr;
	 wire [15:0]execution_unit_0_register_file_0_r9;
	 wire execution_unit_0_register_file_0_n_59_0;
	 wire execution_unit_0_register_file_0_n_59_1;
	 wire execution_unit_0_register_file_0_n_59_2;
	 wire execution_unit_0_register_file_0_n_59_3;
	 wire execution_unit_0_register_file_0_n_59_4;
	 wire execution_unit_0_register_file_0_n_59_5;
	 wire execution_unit_0_register_file_0_n_59_6;
	 wire execution_unit_0_register_file_0_n_59_7;
	 wire execution_unit_0_register_file_0_n_59_8;
	 wire execution_unit_0_register_file_0_n_59_9;
	 wire execution_unit_0_register_file_0_n_59_10;
	 wire execution_unit_0_register_file_0_n_59_11;
	 wire execution_unit_0_register_file_0_n_59_12;
	 wire execution_unit_0_register_file_0_n_59_13;
	 wire execution_unit_0_register_file_0_n_59_14;
	 wire execution_unit_0_register_file_0_n_59_15;
	 wire execution_unit_0_register_file_0_n_59_16;
	 wire execution_unit_0_register_file_0_n_60_0;
	 wire execution_unit_0_register_file_0_n_60_1;
	 wire execution_unit_0_register_file_0_n_62_0;
	 wire execution_unit_0_register_file_0_r10_inc;
	 wire execution_unit_0_register_file_0_r10_wr;
	 wire [15:0]execution_unit_0_register_file_0_r10;
	 wire execution_unit_0_register_file_0_n_66_0;
	 wire execution_unit_0_register_file_0_n_66_1;
	 wire execution_unit_0_register_file_0_n_66_2;
	 wire execution_unit_0_register_file_0_n_66_3;
	 wire execution_unit_0_register_file_0_n_66_4;
	 wire execution_unit_0_register_file_0_n_66_5;
	 wire execution_unit_0_register_file_0_n_66_6;
	 wire execution_unit_0_register_file_0_n_66_7;
	 wire execution_unit_0_register_file_0_n_66_8;
	 wire execution_unit_0_register_file_0_n_66_9;
	 wire execution_unit_0_register_file_0_n_66_10;
	 wire execution_unit_0_register_file_0_n_66_11;
	 wire execution_unit_0_register_file_0_n_66_12;
	 wire execution_unit_0_register_file_0_n_66_13;
	 wire execution_unit_0_register_file_0_n_66_14;
	 wire execution_unit_0_register_file_0_n_66_15;
	 wire execution_unit_0_register_file_0_n_66_16;
	 wire execution_unit_0_register_file_0_n_67_0;
	 wire execution_unit_0_register_file_0_n_67_1;
	 wire execution_unit_0_register_file_0_n_69_0;
	 wire execution_unit_0_register_file_0_r11_inc;
	 wire execution_unit_0_register_file_0_r11_wr;
	 wire [15:0]execution_unit_0_register_file_0_r11;
	 wire execution_unit_0_register_file_0_n_73_0;
	 wire execution_unit_0_register_file_0_n_73_1;
	 wire execution_unit_0_register_file_0_n_73_2;
	 wire execution_unit_0_register_file_0_n_73_3;
	 wire execution_unit_0_register_file_0_n_73_4;
	 wire execution_unit_0_register_file_0_n_73_5;
	 wire execution_unit_0_register_file_0_n_73_6;
	 wire execution_unit_0_register_file_0_n_73_7;
	 wire execution_unit_0_register_file_0_n_73_8;
	 wire execution_unit_0_register_file_0_n_73_9;
	 wire execution_unit_0_register_file_0_n_73_10;
	 wire execution_unit_0_register_file_0_n_73_11;
	 wire execution_unit_0_register_file_0_n_73_12;
	 wire execution_unit_0_register_file_0_n_73_13;
	 wire execution_unit_0_register_file_0_n_73_14;
	 wire execution_unit_0_register_file_0_n_73_15;
	 wire execution_unit_0_register_file_0_n_73_16;
	 wire execution_unit_0_register_file_0_n_74_0;
	 wire execution_unit_0_register_file_0_n_74_1;
	 wire execution_unit_0_register_file_0_n_76_0;
	 wire execution_unit_0_register_file_0_r12_inc;
	 wire execution_unit_0_register_file_0_r12_wr;
	 wire [15:0]execution_unit_0_register_file_0_r12;
	 wire execution_unit_0_register_file_0_n_80_0;
	 wire execution_unit_0_register_file_0_n_80_1;
	 wire execution_unit_0_register_file_0_n_80_2;
	 wire execution_unit_0_register_file_0_n_80_3;
	 wire execution_unit_0_register_file_0_n_80_4;
	 wire execution_unit_0_register_file_0_n_80_5;
	 wire execution_unit_0_register_file_0_n_80_6;
	 wire execution_unit_0_register_file_0_n_80_7;
	 wire execution_unit_0_register_file_0_n_80_8;
	 wire execution_unit_0_register_file_0_n_80_9;
	 wire execution_unit_0_register_file_0_n_80_10;
	 wire execution_unit_0_register_file_0_n_80_11;
	 wire execution_unit_0_register_file_0_n_80_12;
	 wire execution_unit_0_register_file_0_n_80_13;
	 wire execution_unit_0_register_file_0_n_80_14;
	 wire execution_unit_0_register_file_0_n_80_15;
	 wire execution_unit_0_register_file_0_n_80_16;
	 wire execution_unit_0_register_file_0_n_81_0;
	 wire execution_unit_0_register_file_0_n_81_1;
	 wire execution_unit_0_register_file_0_n_83_0;
	 wire execution_unit_0_register_file_0_r13_inc;
	 wire execution_unit_0_register_file_0_r13_wr;
	 wire [15:0]execution_unit_0_register_file_0_r13;
	 wire execution_unit_0_register_file_0_n_87_0;
	 wire execution_unit_0_register_file_0_n_87_1;
	 wire execution_unit_0_register_file_0_n_87_2;
	 wire execution_unit_0_register_file_0_n_87_3;
	 wire execution_unit_0_register_file_0_n_87_4;
	 wire execution_unit_0_register_file_0_n_87_5;
	 wire execution_unit_0_register_file_0_n_87_6;
	 wire execution_unit_0_register_file_0_n_87_7;
	 wire execution_unit_0_register_file_0_n_87_8;
	 wire execution_unit_0_register_file_0_n_87_9;
	 wire execution_unit_0_register_file_0_n_87_10;
	 wire execution_unit_0_register_file_0_n_87_11;
	 wire execution_unit_0_register_file_0_n_87_12;
	 wire execution_unit_0_register_file_0_n_87_13;
	 wire execution_unit_0_register_file_0_n_87_14;
	 wire execution_unit_0_register_file_0_n_87_15;
	 wire execution_unit_0_register_file_0_n_87_16;
	 wire execution_unit_0_register_file_0_n_88_0;
	 wire execution_unit_0_register_file_0_n_88_1;
	 wire execution_unit_0_register_file_0_n_90_0;
	 wire execution_unit_0_register_file_0_r14_inc;
	 wire execution_unit_0_register_file_0_r14_wr;
	 wire [15:0]execution_unit_0_register_file_0_r14;
	 wire execution_unit_0_register_file_0_n_94_0;
	 wire execution_unit_0_register_file_0_n_94_1;
	 wire execution_unit_0_register_file_0_n_94_2;
	 wire execution_unit_0_register_file_0_n_94_3;
	 wire execution_unit_0_register_file_0_n_94_4;
	 wire execution_unit_0_register_file_0_n_94_5;
	 wire execution_unit_0_register_file_0_n_94_6;
	 wire execution_unit_0_register_file_0_n_94_7;
	 wire execution_unit_0_register_file_0_n_94_8;
	 wire execution_unit_0_register_file_0_n_94_9;
	 wire execution_unit_0_register_file_0_n_94_10;
	 wire execution_unit_0_register_file_0_n_94_11;
	 wire execution_unit_0_register_file_0_n_94_12;
	 wire execution_unit_0_register_file_0_n_94_13;
	 wire execution_unit_0_register_file_0_n_94_14;
	 wire execution_unit_0_register_file_0_n_94_15;
	 wire execution_unit_0_register_file_0_n_94_16;
	 wire execution_unit_0_register_file_0_n_95_0;
	 wire execution_unit_0_register_file_0_n_95_1;
	 wire execution_unit_0_register_file_0_n_97_0;
	 wire execution_unit_0_register_file_0_r15_inc;
	 wire execution_unit_0_register_file_0_r15_wr;
	 wire [15:0]execution_unit_0_register_file_0_r15;
	 wire execution_unit_0_register_file_0_n_101_0;
	 wire execution_unit_0_register_file_0_n_101_1;
	 wire execution_unit_0_register_file_0_n_101_2;
	 wire execution_unit_0_register_file_0_n_101_3;
	 wire execution_unit_0_register_file_0_n_101_4;
	 wire execution_unit_0_register_file_0_n_101_5;
	 wire execution_unit_0_register_file_0_n_101_6;
	 wire execution_unit_0_register_file_0_n_101_7;
	 wire execution_unit_0_register_file_0_n_101_8;
	 wire execution_unit_0_register_file_0_n_101_9;
	 wire execution_unit_0_register_file_0_n_101_10;
	 wire execution_unit_0_register_file_0_n_101_11;
	 wire execution_unit_0_register_file_0_n_101_12;
	 wire execution_unit_0_register_file_0_n_101_13;
	 wire execution_unit_0_register_file_0_n_101_14;
	 wire execution_unit_0_register_file_0_n_101_15;
	 wire execution_unit_0_register_file_0_n_101_16;
	 wire execution_unit_0_register_file_0_n_102_0;
	 wire execution_unit_0_register_file_0_n_102_1;
	 wire execution_unit_0_register_file_0_n_104_0;
	 wire execution_unit_0_register_file_0_n_105_0;
	 wire execution_unit_0_register_file_0_n_105_1;
	 wire execution_unit_0_register_file_0_n_105_2;
	 wire execution_unit_0_register_file_0_n_105_3;
	 wire execution_unit_0_register_file_0_n_105_4;
	 wire execution_unit_0_register_file_0_n_105_5;
	 wire execution_unit_0_register_file_0_n_105_6;
	 wire execution_unit_0_register_file_0_n_105_7;
	 wire execution_unit_0_register_file_0_n_105_8;
	 wire execution_unit_0_register_file_0_n_105_9;
	 wire execution_unit_0_register_file_0_n_105_10;
	 wire execution_unit_0_register_file_0_n_105_11;
	 wire execution_unit_0_register_file_0_n_105_12;
	 wire execution_unit_0_register_file_0_n_105_13;
	 wire execution_unit_0_register_file_0_n_105_14;
	 wire execution_unit_0_register_file_0_n_105_15;
	 wire execution_unit_0_register_file_0_n_105_16;
	 wire execution_unit_0_register_file_0_n_105_17;
	 wire execution_unit_0_register_file_0_n_105_18;
	 wire execution_unit_0_register_file_0_n_105_19;
	 wire execution_unit_0_register_file_0_n_105_20;
	 wire execution_unit_0_register_file_0_n_105_21;
	 wire execution_unit_0_register_file_0_n_105_22;
	 wire execution_unit_0_register_file_0_n_105_23;
	 wire execution_unit_0_register_file_0_n_105_24;
	 wire execution_unit_0_register_file_0_n_105_25;
	 wire execution_unit_0_register_file_0_n_105_26;
	 wire execution_unit_0_register_file_0_n_105_27;
	 wire execution_unit_0_register_file_0_n_105_28;
	 wire execution_unit_0_register_file_0_n_105_29;
	 wire execution_unit_0_register_file_0_n_105_30;
	 wire execution_unit_0_register_file_0_n_105_31;
	 wire execution_unit_0_register_file_0_n_105_32;
	 wire execution_unit_0_register_file_0_n_105_33;
	 wire execution_unit_0_register_file_0_n_105_34;
	 wire execution_unit_0_register_file_0_n_105_35;
	 wire execution_unit_0_register_file_0_n_105_36;
	 wire execution_unit_0_register_file_0_n_105_37;
	 wire execution_unit_0_register_file_0_n_105_38;
	 wire execution_unit_0_register_file_0_n_105_39;
	 wire execution_unit_0_register_file_0_n_105_40;
	 wire execution_unit_0_register_file_0_n_105_41;
	 wire execution_unit_0_register_file_0_n_105_42;
	 wire execution_unit_0_register_file_0_n_105_43;
	 wire execution_unit_0_register_file_0_n_105_44;
	 wire execution_unit_0_register_file_0_n_105_45;
	 wire execution_unit_0_register_file_0_n_105_46;
	 wire execution_unit_0_register_file_0_n_105_47;
	 wire execution_unit_0_register_file_0_n_105_48;
	 wire execution_unit_0_register_file_0_n_105_49;
	 wire execution_unit_0_register_file_0_n_105_50;
	 wire execution_unit_0_register_file_0_n_105_51;
	 wire execution_unit_0_register_file_0_n_105_52;
	 wire execution_unit_0_register_file_0_n_105_53;
	 wire execution_unit_0_register_file_0_n_105_54;
	 wire execution_unit_0_register_file_0_n_105_55;
	 wire execution_unit_0_register_file_0_n_105_56;
	 wire execution_unit_0_register_file_0_n_105_57;
	 wire execution_unit_0_register_file_0_n_105_58;
	 wire execution_unit_0_register_file_0_n_105_59;
	 wire execution_unit_0_register_file_0_n_105_60;
	 wire execution_unit_0_register_file_0_n_105_61;
	 wire execution_unit_0_register_file_0_n_105_62;
	 wire execution_unit_0_register_file_0_n_105_63;
	 wire execution_unit_0_register_file_0_n_105_64;
	 wire execution_unit_0_register_file_0_n_105_65;
	 wire execution_unit_0_register_file_0_n_105_66;
	 wire execution_unit_0_register_file_0_n_105_67;
	 wire execution_unit_0_register_file_0_n_105_68;
	 wire execution_unit_0_register_file_0_n_105_69;
	 wire execution_unit_0_register_file_0_n_105_70;
	 wire execution_unit_0_register_file_0_n_105_71;
	 wire execution_unit_0_register_file_0_n_105_72;
	 wire execution_unit_0_register_file_0_n_105_73;
	 wire execution_unit_0_register_file_0_n_105_74;
	 wire execution_unit_0_register_file_0_n_105_75;
	 wire execution_unit_0_register_file_0_n_105_76;
	 wire execution_unit_0_register_file_0_n_105_77;
	 wire execution_unit_0_register_file_0_n_105_78;
	 wire execution_unit_0_register_file_0_n_105_79;
	 wire execution_unit_0_register_file_0_n_105_80;
	 wire execution_unit_0_register_file_0_n_105_81;
	 wire execution_unit_0_register_file_0_n_105_82;
	 wire execution_unit_0_register_file_0_n_105_83;
	 wire execution_unit_0_register_file_0_n_105_84;
	 wire execution_unit_0_register_file_0_n_105_85;
	 wire execution_unit_0_register_file_0_n_105_86;
	 wire execution_unit_0_register_file_0_n_105_87;
	 wire execution_unit_0_register_file_0_n_105_88;
	 wire execution_unit_0_register_file_0_n_105_89;
	 wire execution_unit_0_register_file_0_n_105_90;
	 wire execution_unit_0_register_file_0_n_105_91;
	 wire execution_unit_0_register_file_0_n_105_92;
	 wire execution_unit_0_register_file_0_n_105_93;
	 wire execution_unit_0_register_file_0_n_105_94;
	 wire execution_unit_0_register_file_0_n_105_95;
	 wire execution_unit_0_register_file_0_n_105_96;
	 wire execution_unit_0_register_file_0_n_105_97;
	 wire execution_unit_0_register_file_0_n_105_98;
	 wire execution_unit_0_register_file_0_n_105_99;
	 wire execution_unit_0_register_file_0_n_105_100;
	 wire execution_unit_0_register_file_0_n_105_101;
	 wire execution_unit_0_register_file_0_n_105_102;
	 wire execution_unit_0_register_file_0_n_105_103;
	 wire execution_unit_0_register_file_0_n_105_104;
	 wire execution_unit_0_register_file_0_n_105_105;
	 wire execution_unit_0_register_file_0_n_105_106;
	 wire execution_unit_0_register_file_0_n_105_107;
	 wire execution_unit_0_register_file_0_n_105_108;
	 wire execution_unit_0_register_file_0_n_105_109;
	 wire execution_unit_0_register_file_0_n_105_110;
	 wire execution_unit_0_register_file_0_n_105_111;
	 wire execution_unit_0_register_file_0_n_105_112;
	 wire execution_unit_0_register_file_0_n_105_113;
	 wire execution_unit_0_register_file_0_n_105_114;
	 wire execution_unit_0_register_file_0_n_105_115;
	 wire execution_unit_0_register_file_0_n_105_116;
	 wire execution_unit_0_register_file_0_n_105_117;
	 wire execution_unit_0_register_file_0_n_105_118;
	 wire execution_unit_0_register_file_0_n_105_119;
	 wire execution_unit_0_register_file_0_n_105_120;
	 wire execution_unit_0_register_file_0_n_105_121;
	 wire execution_unit_0_register_file_0_n_105_122;
	 wire execution_unit_0_register_file_0_n_105_123;
	 wire execution_unit_0_register_file_0_n_105_124;
	 wire execution_unit_0_register_file_0_n_105_125;
	 wire execution_unit_0_register_file_0_n_105_126;
	 wire execution_unit_0_register_file_0_n_105_127;
	 wire execution_unit_0_register_file_0_n_105_128;
	 wire execution_unit_0_register_file_0_n_105_129;
	 wire execution_unit_0_register_file_0_n_105_130;
	 wire execution_unit_0_register_file_0_n_105_131;
	 wire execution_unit_0_register_file_0_n_105_132;
	 wire execution_unit_0_register_file_0_n_105_133;
	 wire execution_unit_0_register_file_0_n_105_134;
	 wire execution_unit_0_register_file_0_n_105_135;
	 wire execution_unit_0_register_file_0_n_105_136;
	 wire execution_unit_0_register_file_0_n_105_137;
	 wire execution_unit_0_register_file_0_n_105_138;
	 wire execution_unit_0_register_file_0_n_105_139;
	 wire execution_unit_0_register_file_0_n_105_140;
	 wire execution_unit_0_register_file_0_n_105_141;
	 wire execution_unit_0_register_file_0_n_105_142;
	 wire execution_unit_0_register_file_0_n_105_143;
	 wire execution_unit_0_register_file_0_n_105_144;
	 wire execution_unit_0_register_file_0_n_105_145;
	 wire execution_unit_0_register_file_0_n_105_146;
	 wire execution_unit_0_register_file_0_n_105_147;
	 wire execution_unit_0_register_file_0_n_105_148;
	 wire execution_unit_0_register_file_0_n_105_149;
	 wire execution_unit_0_register_file_0_n_105_150;
	 wire execution_unit_0_register_file_0_n_105_151;
	 wire execution_unit_0_register_file_0_n_105_152;
	 wire execution_unit_0_register_file_0_n_105_153;
	 wire execution_unit_0_register_file_0_n_105_154;
	 wire execution_unit_0_register_file_0_n_105_155;
	 wire execution_unit_0_register_file_0_n_105_156;
	 wire execution_unit_0_register_file_0_n_105_157;
	 wire execution_unit_0_register_file_0_n_105_158;
	 wire execution_unit_0_register_file_0_n_105_159;
	 wire execution_unit_0_register_file_0_n_105_160;
	 wire execution_unit_0_register_file_0_n_105_161;
	 wire execution_unit_0_register_file_0_n_105_162;
	 wire execution_unit_0_register_file_0_n_105_163;
	 wire execution_unit_0_register_file_0_n_105_164;
	 wire execution_unit_0_register_file_0_n_105_165;
	 wire execution_unit_0_register_file_0_n_105_166;
	 wire execution_unit_0_register_file_0_n_105_167;
	 wire execution_unit_0_register_file_0_n_105_168;
	 wire execution_unit_0_register_file_0_n_105_169;
	 wire execution_unit_0_register_file_0_n_105_170;
	 wire execution_unit_0_register_file_0_n_105_171;
	 wire execution_unit_0_register_file_0_n_105_172;
	 wire execution_unit_0_register_file_0_n_105_173;
	 wire execution_unit_0_register_file_0_n_105_174;
	 wire execution_unit_0_register_file_0_n_105_175;
	 wire execution_unit_0_register_file_0_n_105_176;
	 wire execution_unit_0_register_file_0_n_105_177;
	 wire execution_unit_0_register_file_0_n_105_178;
	 wire execution_unit_0_register_file_0_n_105_179;
	 wire execution_unit_0_register_file_0_n_105_180;
	 wire execution_unit_0_register_file_0_n_105_181;
	 wire execution_unit_0_register_file_0_n_105_182;
	 wire execution_unit_0_register_file_0_n_105_183;
	 wire execution_unit_0_register_file_0_n_105_184;
	 wire execution_unit_0_register_file_0_n_105_185;
	 wire execution_unit_0_register_file_0_n_105_186;
	 wire execution_unit_0_register_file_0_n_105_187;
	 wire execution_unit_0_register_file_0_n_105_188;
	 wire execution_unit_0_register_file_0_n_105_189;
	 wire execution_unit_0_register_file_0_n_105_190;
	 wire execution_unit_0_register_file_0_n_105_191;
	 wire execution_unit_0_register_file_0_n_105_192;
	 wire execution_unit_0_register_file_0_n_105_193;
	 wire execution_unit_0_register_file_0_n_105_194;
	 wire execution_unit_0_register_file_0_n_105_195;
	 wire execution_unit_0_register_file_0_n_105_196;
	 wire execution_unit_0_register_file_0_n_105_197;
	 wire execution_unit_0_register_file_0_n_105_198;
	 wire execution_unit_0_register_file_0_n_105_199;
	 wire execution_unit_0_register_file_0_n_105_200;
	 wire execution_unit_0_register_file_0_n_105_201;
	 wire execution_unit_0_register_file_0_n_105_202;
	 wire execution_unit_0_register_file_0_n_105_203;
	 wire execution_unit_0_register_file_0_n_105_204;
	 wire execution_unit_0_register_file_0_n_105_205;
	 wire execution_unit_0_register_file_0_n_105_206;
	 wire execution_unit_0_register_file_0_n_105_207;
	 wire execution_unit_0_register_file_0_n_105_208;
	 wire execution_unit_0_register_file_0_n_105_209;
	 wire execution_unit_0_register_file_0_n_105_210;
	 wire execution_unit_0_register_file_0_n_105_211;
	 wire execution_unit_0_register_file_0_n_105_212;
	 wire execution_unit_0_register_file_0_n_105_213;
	 wire execution_unit_0_register_file_0_n_105_214;
	 wire execution_unit_0_register_file_0_n_105_215;
	 wire execution_unit_0_register_file_0_n_105_216;
	 wire execution_unit_0_register_file_0_n_105_217;
	 wire execution_unit_0_register_file_0_n_105_218;
	 wire execution_unit_0_register_file_0_n_105_219;
	 wire execution_unit_0_register_file_0_n_105_220;
	 wire execution_unit_0_register_file_0_n_105_221;
	 wire execution_unit_0_register_file_0_n_105_222;
	 wire execution_unit_0_register_file_0_n_105_223;
	 wire execution_unit_0_register_file_0_n_105_224;
	 wire execution_unit_0_register_file_0_n_105_225;
	 wire execution_unit_0_register_file_0_n_105_226;
	 wire execution_unit_0_register_file_0_n_105_227;
	 wire execution_unit_0_register_file_0_n_105_228;
	 wire execution_unit_0_register_file_0_n_105_229;
	 wire execution_unit_0_register_file_0_n_105_230;
	 wire execution_unit_0_register_file_0_n_105_231;
	 wire execution_unit_0_register_file_0_n_105_232;
	 wire execution_unit_0_register_file_0_n_105_233;
	 wire execution_unit_0_register_file_0_n_105_234;
	 wire execution_unit_0_register_file_0_n_105_235;
	 wire execution_unit_0_register_file_0_n_105_236;
	 wire execution_unit_0_register_file_0_n_105_237;
	 wire execution_unit_0_register_file_0_n_105_238;
	 wire execution_unit_0_register_file_0_n_105_239;
	 wire execution_unit_0_register_file_0_n_105_240;
	 wire execution_unit_0_register_file_0_n_105_241;
	 wire execution_unit_0_register_file_0_n_105_242;
	 wire execution_unit_0_register_file_0_n_105_243;
	 wire execution_unit_0_register_file_0_n_105_244;
	 wire execution_unit_0_register_file_0_n_105_245;
	 wire execution_unit_0_register_file_0_n_105_246;
	 wire execution_unit_0_register_file_0_n_105_247;
	 wire execution_unit_0_register_file_0_n_105_248;
	 wire execution_unit_0_register_file_0_n_105_249;
	 wire execution_unit_0_register_file_0_n_105_250;
	 wire execution_unit_0_register_file_0_n_105_251;
	 wire execution_unit_0_register_file_0_n_105_252;
	 wire execution_unit_0_register_file_0_n_105_253;
	 wire execution_unit_0_register_file_0_n_105_254;
	 wire execution_unit_0_register_file_0_n_105_255;
	 wire execution_unit_0_register_file_0_n_105_256;
	 wire execution_unit_0_register_file_0_n_105_257;
	 wire execution_unit_0_register_file_0_n_105_258;
	 wire execution_unit_0_register_file_0_n_105_259;
	 wire execution_unit_0_register_file_0_n_105_260;
	 wire execution_unit_0_register_file_0_n_105_261;
	 wire execution_unit_0_register_file_0_n_105_262;
	 wire execution_unit_0_register_file_0_n_105_263;
	 wire execution_unit_0_register_file_0_n_105_264;
	 wire execution_unit_0_register_file_0_n_105_265;
	 wire execution_unit_0_register_file_0_n_105_266;
	 wire execution_unit_0_register_file_0_n_105_267;
	 wire execution_unit_0_register_file_0_n_105_268;
	 wire execution_unit_0_register_file_0_n_105_269;
	 wire execution_unit_0_register_file_0_n_105_270;
	 wire execution_unit_0_register_file_0_n_105_271;
	 wire execution_unit_0_register_file_0_n_105_272;
	 wire execution_unit_0_register_file_0_n_105_273;
	 wire execution_unit_0_register_file_0_n_105_274;
	 wire execution_unit_0_register_file_0_n_105_275;
	 wire execution_unit_0_register_file_0_n_105_276;
	 wire execution_unit_0_register_file_0_n_105_277;
	 wire execution_unit_0_register_file_0_n_105_278;
	 wire execution_unit_0_register_file_0_n_105_279;
	 wire execution_unit_0_register_file_0_n_105_280;
	 wire execution_unit_0_register_file_0_n_105_281;
	 wire execution_unit_0_register_file_0_n_105_282;
	 wire execution_unit_0_register_file_0_n_105_283;
	 wire execution_unit_0_register_file_0_n_105_284;
	 wire execution_unit_0_register_file_0_n_105_285;
	 wire execution_unit_0_register_file_0_n_105_286;
	 wire execution_unit_0_register_file_0_n_105_287;
	 wire execution_unit_0_register_file_0_n_105_288;
	 wire execution_unit_0_register_file_0_n_105_289;
	 wire execution_unit_0_register_file_0_n_105_290;
	 wire execution_unit_0_register_file_0_n_105_291;
	 wire execution_unit_0_register_file_0_n_105_292;
	 wire execution_unit_0_register_file_0_n_105_293;
	 wire execution_unit_0_register_file_0_n_105_294;
	 wire execution_unit_0_register_file_0_n_105_295;
	 wire execution_unit_0_register_file_0_n_105_296;
	 wire execution_unit_0_register_file_0_n_105_297;
	 wire execution_unit_0_register_file_0_n_105_298;
	 wire execution_unit_0_register_file_0_n_105_299;
	 wire execution_unit_0_register_file_0_n_105_300;
	 wire execution_unit_0_register_file_0_n_105_301;
	 wire execution_unit_0_register_file_0_n_105_302;
	 wire execution_unit_0_register_file_0_n_105_303;
	 wire execution_unit_0_register_file_0_n_105_304;
	 wire execution_unit_0_register_file_0_n_105_305;
	 wire execution_unit_0_register_file_0_n_105_306;
	 wire execution_unit_0_register_file_0_n_105_307;
	 wire execution_unit_0_register_file_0_n_105_308;
	 wire execution_unit_0_register_file_0_n_105_309;
	 wire execution_unit_0_register_file_0_n_105_310;
	 wire execution_unit_0_register_file_0_n_105_311;
	 wire execution_unit_0_register_file_0_n_105_312;
	 wire execution_unit_0_register_file_0_n_105_313;
	 wire execution_unit_0_register_file_0_n_105_314;
	 wire execution_unit_0_register_file_0_n_105_315;
	 wire execution_unit_0_register_file_0_n_105_316;
	 wire execution_unit_0_register_file_0_n_105_317;
	 wire execution_unit_0_register_file_0_n_105_318;
	 wire execution_unit_0_register_file_0_n_105_319;
	 wire execution_unit_0_register_file_0_n_106_0;
	 wire execution_unit_0_register_file_0_n_106_1;
	 wire execution_unit_0_register_file_0_n_106_2;
	 wire execution_unit_0_register_file_0_n_106_3;
	 wire execution_unit_0_register_file_0_n_106_4;
	 wire execution_unit_0_register_file_0_n_106_5;
	 wire execution_unit_0_register_file_0_n_106_6;
	 wire execution_unit_0_register_file_0_n_106_7;
	 wire execution_unit_0_register_file_0_n_106_8;
	 wire execution_unit_0_register_file_0_n_106_9;
	 wire execution_unit_0_register_file_0_n_106_10;
	 wire execution_unit_0_register_file_0_n_106_11;
	 wire execution_unit_0_register_file_0_n_106_12;
	 wire execution_unit_0_register_file_0_n_106_13;
	 wire [15:0]execution_unit_0_register_file_0_r1;
	 wire execution_unit_0_register_file_0_n_108_0;
	 wire execution_unit_0_register_file_0_n_109_0;
	 wire execution_unit_0_register_file_0_n_109_1;
	 wire execution_unit_0_register_file_0_n_109_2;
	 wire execution_unit_0_register_file_0_n_109_3;
	 wire execution_unit_0_register_file_0_n_109_4;
	 wire execution_unit_0_register_file_0_n_109_5;
	 wire execution_unit_0_register_file_0_n_109_6;
	 wire execution_unit_0_register_file_0_n_109_7;
	 wire execution_unit_0_register_file_0_n_109_8;
	 wire execution_unit_0_register_file_0_n_109_9;
	 wire execution_unit_0_register_file_0_n_109_10;
	 wire execution_unit_0_register_file_0_n_109_11;
	 wire execution_unit_0_register_file_0_n_109_12;
	 wire execution_unit_0_register_file_0_n_109_13;
	 wire execution_unit_0_register_file_0_n_109_14;
	 wire execution_unit_0_register_file_0_n_110_0;
	 wire execution_unit_0_register_file_0_n_110_1;
	 wire execution_unit_0_register_file_0_n_110_2;
	 wire execution_unit_0_register_file_0_n_112_0;
	 wire execution_unit_0_register_file_0_n_112_1;
	 wire execution_unit_0_register_file_0_n_112_2;
	 wire execution_unit_0_register_file_0_n_112_3;
	 wire execution_unit_0_register_file_0_n_112_4;
	 wire execution_unit_0_register_file_0_n_112_5;
	 wire execution_unit_0_register_file_0_n_112_6;
	 wire execution_unit_0_register_file_0_n_112_7;
	 wire execution_unit_0_register_file_0_n_112_8;
	 wire execution_unit_0_register_file_0_n_112_9;
	 wire execution_unit_0_register_file_0_n_112_10;
	 wire execution_unit_0_register_file_0_n_112_11;
	 wire execution_unit_0_register_file_0_n_112_12;
	 wire execution_unit_0_register_file_0_n_112_13;
	 wire execution_unit_0_register_file_0_n_112_14;
	 wire execution_unit_0_register_file_0_n_112_15;
	 wire execution_unit_0_register_file_0_n_112_16;
	 wire execution_unit_0_register_file_0_n_112_17;
	 wire execution_unit_0_register_file_0_n_112_18;
	 wire execution_unit_0_register_file_0_n_112_19;
	 wire execution_unit_0_register_file_0_n_112_20;
	 wire execution_unit_0_register_file_0_n_112_21;
	 wire execution_unit_0_register_file_0_n_112_22;
	 wire execution_unit_0_register_file_0_n_112_23;
	 wire execution_unit_0_register_file_0_n_112_24;
	 wire execution_unit_0_register_file_0_n_112_25;
	 wire execution_unit_0_register_file_0_n_112_26;
	 wire execution_unit_0_register_file_0_n_112_27;
	 wire execution_unit_0_register_file_0_n_112_28;
	 wire execution_unit_0_register_file_0_n_112_29;
	 wire execution_unit_0_register_file_0_n_112_30;
	 wire execution_unit_0_register_file_0_n_112_31;
	 wire execution_unit_0_register_file_0_n_112_32;
	 wire execution_unit_0_register_file_0_n_112_33;
	 wire execution_unit_0_register_file_0_n_112_34;
	 wire execution_unit_0_register_file_0_n_112_35;
	 wire execution_unit_0_register_file_0_n_112_36;
	 wire execution_unit_0_register_file_0_n_112_37;
	 wire execution_unit_0_register_file_0_n_112_38;
	 wire execution_unit_0_register_file_0_n_112_39;
	 wire execution_unit_0_register_file_0_n_112_40;
	 wire execution_unit_0_register_file_0_n_112_41;
	 wire execution_unit_0_register_file_0_n_112_42;
	 wire execution_unit_0_register_file_0_n_112_43;
	 wire execution_unit_0_register_file_0_n_112_44;
	 wire execution_unit_0_register_file_0_n_112_45;
	 wire execution_unit_0_register_file_0_n_112_46;
	 wire execution_unit_0_register_file_0_n_112_47;
	 wire execution_unit_0_register_file_0_n_112_48;
	 wire execution_unit_0_register_file_0_n_112_49;
	 wire execution_unit_0_register_file_0_n_112_50;
	 wire execution_unit_0_register_file_0_n_112_51;
	 wire execution_unit_0_register_file_0_n_112_52;
	 wire execution_unit_0_register_file_0_n_112_53;
	 wire execution_unit_0_register_file_0_n_112_54;
	 wire execution_unit_0_register_file_0_n_112_55;
	 wire execution_unit_0_register_file_0_n_112_56;
	 wire execution_unit_0_register_file_0_n_112_57;
	 wire execution_unit_0_register_file_0_n_112_58;
	 wire execution_unit_0_register_file_0_n_112_59;
	 wire execution_unit_0_register_file_0_n_112_60;
	 wire execution_unit_0_register_file_0_n_112_61;
	 wire execution_unit_0_register_file_0_n_112_62;
	 wire execution_unit_0_register_file_0_n_112_63;
	 wire execution_unit_0_register_file_0_n_112_64;
	 wire execution_unit_0_register_file_0_n_112_65;
	 wire execution_unit_0_register_file_0_n_112_66;
	 wire execution_unit_0_register_file_0_n_112_67;
	 wire execution_unit_0_register_file_0_n_112_68;
	 wire execution_unit_0_register_file_0_n_112_69;
	 wire execution_unit_0_register_file_0_n_112_70;
	 wire execution_unit_0_register_file_0_n_112_71;
	 wire execution_unit_0_register_file_0_n_112_72;
	 wire execution_unit_0_register_file_0_n_112_73;
	 wire execution_unit_0_register_file_0_n_112_74;
	 wire execution_unit_0_register_file_0_n_112_75;
	 wire execution_unit_0_register_file_0_n_112_76;
	 wire execution_unit_0_register_file_0_n_112_77;
	 wire execution_unit_0_register_file_0_n_112_78;
	 wire execution_unit_0_register_file_0_n_112_79;
	 wire execution_unit_0_register_file_0_n_112_80;
	 wire execution_unit_0_register_file_0_n_112_81;
	 wire execution_unit_0_register_file_0_n_112_82;
	 wire execution_unit_0_register_file_0_n_112_83;
	 wire execution_unit_0_register_file_0_n_112_84;
	 wire execution_unit_0_register_file_0_n_112_85;
	 wire execution_unit_0_register_file_0_n_112_86;
	 wire execution_unit_0_register_file_0_n_112_87;
	 wire execution_unit_0_register_file_0_n_112_88;
	 wire execution_unit_0_register_file_0_n_112_89;
	 wire execution_unit_0_register_file_0_n_112_90;
	 wire execution_unit_0_register_file_0_n_112_91;
	 wire execution_unit_0_register_file_0_n_112_92;
	 wire execution_unit_0_register_file_0_n_112_93;
	 wire execution_unit_0_register_file_0_n_112_94;
	 wire execution_unit_0_register_file_0_n_112_95;
	 wire execution_unit_0_register_file_0_n_112_96;
	 wire execution_unit_0_register_file_0_n_112_97;
	 wire execution_unit_0_register_file_0_n_112_98;
	 wire execution_unit_0_register_file_0_n_112_99;
	 wire execution_unit_0_register_file_0_n_112_100;
	 wire execution_unit_0_register_file_0_n_112_101;
	 wire execution_unit_0_register_file_0_n_112_102;
	 wire execution_unit_0_register_file_0_n_112_103;
	 wire execution_unit_0_register_file_0_n_112_104;
	 wire execution_unit_0_register_file_0_n_112_105;
	 wire execution_unit_0_register_file_0_n_112_106;
	 wire execution_unit_0_register_file_0_n_112_107;
	 wire execution_unit_0_register_file_0_n_112_108;
	 wire execution_unit_0_register_file_0_n_112_109;
	 wire execution_unit_0_register_file_0_n_112_110;
	 wire execution_unit_0_register_file_0_n_112_111;
	 wire execution_unit_0_register_file_0_n_112_112;
	 wire execution_unit_0_register_file_0_n_112_113;
	 wire execution_unit_0_register_file_0_n_112_114;
	 wire execution_unit_0_register_file_0_n_112_115;
	 wire execution_unit_0_register_file_0_n_112_116;
	 wire execution_unit_0_register_file_0_n_112_117;
	 wire execution_unit_0_register_file_0_n_112_118;
	 wire execution_unit_0_register_file_0_n_112_119;
	 wire execution_unit_0_register_file_0_n_112_120;
	 wire execution_unit_0_register_file_0_n_112_121;
	 wire execution_unit_0_register_file_0_n_112_122;
	 wire execution_unit_0_register_file_0_n_112_123;
	 wire execution_unit_0_register_file_0_n_112_124;
	 wire execution_unit_0_register_file_0_n_112_125;
	 wire execution_unit_0_register_file_0_n_112_126;
	 wire execution_unit_0_register_file_0_n_112_127;
	 wire execution_unit_0_register_file_0_n_112_128;
	 wire execution_unit_0_register_file_0_n_112_129;
	 wire execution_unit_0_register_file_0_n_112_130;
	 wire execution_unit_0_register_file_0_n_112_131;
	 wire execution_unit_0_register_file_0_n_112_132;
	 wire execution_unit_0_register_file_0_n_112_133;
	 wire execution_unit_0_register_file_0_n_112_134;
	 wire execution_unit_0_register_file_0_n_112_135;
	 wire execution_unit_0_register_file_0_n_112_136;
	 wire execution_unit_0_register_file_0_n_112_137;
	 wire execution_unit_0_register_file_0_n_112_138;
	 wire execution_unit_0_register_file_0_n_112_139;
	 wire execution_unit_0_register_file_0_n_112_140;
	 wire execution_unit_0_register_file_0_n_112_141;
	 wire execution_unit_0_register_file_0_n_112_142;
	 wire execution_unit_0_register_file_0_n_112_143;
	 wire execution_unit_0_register_file_0_n_112_144;
	 wire execution_unit_0_register_file_0_n_112_145;
	 wire execution_unit_0_register_file_0_n_112_146;
	 wire execution_unit_0_register_file_0_n_112_147;
	 wire execution_unit_0_register_file_0_n_112_148;
	 wire execution_unit_0_register_file_0_n_112_149;
	 wire execution_unit_0_register_file_0_n_112_150;
	 wire execution_unit_0_register_file_0_n_112_151;
	 wire execution_unit_0_register_file_0_n_112_152;
	 wire execution_unit_0_register_file_0_n_112_153;
	 wire execution_unit_0_register_file_0_n_112_154;
	 wire execution_unit_0_register_file_0_n_112_155;
	 wire execution_unit_0_register_file_0_n_112_156;
	 wire execution_unit_0_register_file_0_n_112_157;
	 wire execution_unit_0_register_file_0_n_112_158;
	 wire execution_unit_0_register_file_0_n_112_159;
	 wire execution_unit_0_register_file_0_n_112_160;
	 wire execution_unit_0_register_file_0_n_112_161;
	 wire execution_unit_0_register_file_0_n_112_162;
	 wire execution_unit_0_register_file_0_n_112_163;
	 wire execution_unit_0_register_file_0_n_112_164;
	 wire execution_unit_0_register_file_0_n_112_165;
	 wire execution_unit_0_register_file_0_n_112_166;
	 wire execution_unit_0_register_file_0_n_112_167;
	 wire execution_unit_0_register_file_0_n_112_168;
	 wire execution_unit_0_register_file_0_n_112_169;
	 wire execution_unit_0_register_file_0_n_112_170;
	 wire execution_unit_0_register_file_0_n_112_171;
	 wire execution_unit_0_register_file_0_n_112_172;
	 wire execution_unit_0_register_file_0_n_112_173;
	 wire execution_unit_0_register_file_0_n_112_174;
	 wire execution_unit_0_register_file_0_n_112_175;
	 wire execution_unit_0_register_file_0_n_112_176;
	 wire execution_unit_0_register_file_0_n_112_177;
	 wire execution_unit_0_register_file_0_n_112_178;
	 wire execution_unit_0_register_file_0_n_112_179;
	 wire execution_unit_0_register_file_0_n_112_180;
	 wire execution_unit_0_register_file_0_n_112_181;
	 wire execution_unit_0_register_file_0_n_112_182;
	 wire execution_unit_0_register_file_0_n_112_183;
	 wire execution_unit_0_register_file_0_n_112_184;
	 wire execution_unit_0_register_file_0_n_112_185;
	 wire execution_unit_0_register_file_0_n_112_186;
	 wire execution_unit_0_register_file_0_n_112_187;
	 wire execution_unit_0_register_file_0_n_112_188;
	 wire execution_unit_0_register_file_0_n_112_189;
	 wire execution_unit_0_register_file_0_n_112_190;
	 wire execution_unit_0_register_file_0_n_112_191;
	 wire execution_unit_0_register_file_0_n_112_192;
	 wire execution_unit_0_register_file_0_n_112_193;
	 wire execution_unit_0_register_file_0_n_112_194;
	 wire execution_unit_0_register_file_0_n_112_195;
	 wire execution_unit_0_register_file_0_n_112_196;
	 wire execution_unit_0_register_file_0_n_112_197;
	 wire execution_unit_0_register_file_0_n_112_198;
	 wire execution_unit_0_register_file_0_n_112_199;
	 wire execution_unit_0_register_file_0_n_112_200;
	 wire execution_unit_0_register_file_0_n_112_201;
	 wire execution_unit_0_register_file_0_n_112_202;
	 wire execution_unit_0_register_file_0_n_112_203;
	 wire execution_unit_0_register_file_0_n_112_204;
	 wire execution_unit_0_register_file_0_n_112_205;
	 wire execution_unit_0_register_file_0_n_112_206;
	 wire execution_unit_0_register_file_0_n_112_207;
	 wire execution_unit_0_register_file_0_n_112_208;
	 wire execution_unit_0_register_file_0_n_112_209;
	 wire execution_unit_0_register_file_0_n_112_210;
	 wire execution_unit_0_register_file_0_n_112_211;
	 wire execution_unit_0_register_file_0_n_112_212;
	 wire execution_unit_0_register_file_0_n_112_213;
	 wire execution_unit_0_register_file_0_n_112_214;
	 wire execution_unit_0_register_file_0_n_112_215;
	 wire execution_unit_0_register_file_0_n_112_216;
	 wire execution_unit_0_register_file_0_n_112_217;
	 wire execution_unit_0_register_file_0_n_112_218;
	 wire execution_unit_0_register_file_0_n_112_219;
	 wire execution_unit_0_register_file_0_n_112_220;
	 wire execution_unit_0_register_file_0_n_112_221;
	 wire execution_unit_0_register_file_0_n_112_222;
	 wire execution_unit_0_register_file_0_n_112_223;
	 wire execution_unit_0_register_file_0_n_112_224;
	 wire execution_unit_0_register_file_0_n_112_225;
	 wire execution_unit_0_register_file_0_n_112_226;
	 wire execution_unit_0_register_file_0_n_112_227;
	 wire execution_unit_0_register_file_0_n_112_228;
	 wire execution_unit_0_register_file_0_n_112_229;
	 wire execution_unit_0_register_file_0_n_112_230;
	 wire execution_unit_0_register_file_0_n_112_231;
	 wire execution_unit_0_register_file_0_n_112_232;
	 wire execution_unit_0_register_file_0_n_112_233;
	 wire execution_unit_0_register_file_0_n_112_234;
	 wire execution_unit_0_register_file_0_n_112_235;
	 wire execution_unit_0_register_file_0_n_112_236;
	 wire execution_unit_0_register_file_0_n_112_237;
	 wire execution_unit_0_register_file_0_n_112_238;
	 wire execution_unit_0_register_file_0_n_112_239;
	 wire execution_unit_0_register_file_0_n_112_240;
	 wire execution_unit_0_register_file_0_n_112_241;
	 wire execution_unit_0_register_file_0_n_112_242;
	 wire execution_unit_0_register_file_0_n_112_243;
	 wire execution_unit_0_register_file_0_n_112_244;
	 wire execution_unit_0_register_file_0_n_112_245;
	 wire execution_unit_0_register_file_0_n_112_246;
	 wire execution_unit_0_register_file_0_n_112_247;
	 wire execution_unit_0_register_file_0_n_112_248;
	 wire execution_unit_0_register_file_0_n_112_249;
	 wire execution_unit_0_register_file_0_n_112_250;
	 wire execution_unit_0_register_file_0_n_112_251;
	 wire execution_unit_0_register_file_0_n_112_252;
	 wire execution_unit_0_register_file_0_n_112_253;
	 wire execution_unit_0_register_file_0_n_112_254;
	 wire execution_unit_0_register_file_0_n_112_255;
	 wire execution_unit_0_register_file_0_n_112_256;
	 wire execution_unit_0_register_file_0_n_112_257;
	 wire execution_unit_0_register_file_0_n_112_258;
	 wire execution_unit_0_register_file_0_n_112_259;
	 wire execution_unit_0_register_file_0_n_112_260;
	 wire execution_unit_0_register_file_0_n_112_261;
	 wire execution_unit_0_register_file_0_n_112_262;
	 wire execution_unit_0_register_file_0_n_112_263;
	 wire execution_unit_0_register_file_0_n_112_264;
	 wire execution_unit_0_register_file_0_n_112_265;
	 wire execution_unit_0_register_file_0_n_112_266;
	 wire execution_unit_0_register_file_0_n_112_267;
	 wire execution_unit_0_register_file_0_n_112_268;
	 wire execution_unit_0_register_file_0_n_112_269;
	 wire execution_unit_0_register_file_0_n_112_270;
	 wire execution_unit_0_register_file_0_n_112_271;
	 wire execution_unit_0_register_file_0_n_112_272;
	 wire execution_unit_0_register_file_0_n_112_273;
	 wire execution_unit_0_register_file_0_n_112_274;
	 wire execution_unit_0_register_file_0_n_112_275;
	 wire execution_unit_0_register_file_0_n_112_276;
	 wire execution_unit_0_register_file_0_n_112_277;
	 wire execution_unit_0_register_file_0_n_112_278;
	 wire execution_unit_0_register_file_0_n_112_279;
	 wire execution_unit_0_register_file_0_n_112_280;
	 wire execution_unit_0_register_file_0_n_112_281;
	 wire execution_unit_0_register_file_0_n_112_282;
	 wire execution_unit_0_register_file_0_n_112_283;
	 wire execution_unit_0_register_file_0_n_112_284;
	 wire execution_unit_0_register_file_0_n_112_285;
	 wire execution_unit_0_register_file_0_n_112_286;
	 wire execution_unit_0_register_file_0_n_112_287;
	 wire execution_unit_0_register_file_0_n_112_288;
	 wire execution_unit_0_register_file_0_n_112_289;
	 wire execution_unit_0_register_file_0_n_112_290;
	 wire execution_unit_0_register_file_0_n_112_291;
	 wire execution_unit_0_register_file_0_n_112_292;
	 wire execution_unit_0_register_file_0_n_112_293;
	 wire execution_unit_0_register_file_0_n_112_294;
	 wire execution_unit_0_register_file_0_n_112_295;
	 wire execution_unit_0_register_file_0_n_112_296;
	 wire execution_unit_0_register_file_0_n_112_297;
	 wire execution_unit_0_register_file_0_n_112_298;
	 wire execution_unit_0_register_file_0_n_112_299;
	 wire execution_unit_0_register_file_0_n_112_300;
	 wire execution_unit_0_register_file_0_n_112_301;
	 wire execution_unit_0_register_file_0_n_112_302;
	 wire execution_unit_0_register_file_0_n_112_303;
	 wire execution_unit_0_register_file_0_n_112_304;
	 wire execution_unit_0_register_file_0_n_112_305;
	 wire execution_unit_0_register_file_0_n_112_306;
	 wire execution_unit_0_register_file_0_n_112_307;
	 wire execution_unit_0_register_file_0_n_112_308;
	 wire execution_unit_0_register_file_0_n_112_309;
	 wire execution_unit_0_register_file_0_n_112_310;
	 wire execution_unit_0_register_file_0_n_112_311;
	 wire execution_unit_0_register_file_0_n_112_312;
	 wire execution_unit_0_register_file_0_n_112_313;
	 wire execution_unit_0_register_file_0_n_112_314;
	 wire execution_unit_0_register_file_0_n_112_315;
	 wire execution_unit_0_register_file_0_n_112_316;
	 wire execution_unit_0_register_file_0_n_112_317;
	 wire execution_unit_0_register_file_0_n_112_318;
	 wire execution_unit_0_register_file_0_n_112_319;
	 wire execution_unit_0_register_file_0_n_7;
	 wire execution_unit_0_register_file_0_n_17;
	 wire execution_unit_0_register_file_0_n_8;
	 wire execution_unit_0_register_file_0_n_16;
	 wire execution_unit_0_register_file_0_n_24;
	 wire execution_unit_0_register_file_0_n_22;
	 wire execution_unit_0_register_file_0_n_23;
	 wire execution_unit_0_register_file_0_n_21;
	 wire execution_unit_0_register_file_0_n_0;
	 wire execution_unit_0_register_file_0_n_272;
	 wire execution_unit_0_register_file_0_n_271;
	 wire execution_unit_0_register_file_0_n_41;
	 wire execution_unit_0_register_file_0_n_44;
	 wire execution_unit_0_register_file_0_n_27;
	 wire execution_unit_0_register_file_0_n_2;
	 wire execution_unit_0_register_file_0_n_39;
	 wire execution_unit_0_register_file_0_n_4;
	 wire execution_unit_0_register_file_0_n_37;
	 wire execution_unit_0_register_file_0_n_6;
	 wire execution_unit_0_register_file_0_n_35;
	 wire execution_unit_0_register_file_0_n_19;
	 wire execution_unit_0_register_file_0_n_33;
	 wire execution_unit_0_register_file_0_n_31;
	 wire execution_unit_0_register_file_0_n_25;
	 wire execution_unit_0_register_file_0_n_26;
	 wire execution_unit_0_register_file_0_n_29;
	 wire execution_unit_0_register_file_0_n_10;
	 wire execution_unit_0_register_file_0_n_14;
	 wire execution_unit_0_register_file_0_n_255;
	 wire execution_unit_0_register_file_0_n_273;
	 wire execution_unit_0_register_file_0_n_288;
	 wire execution_unit_0_register_file_0_n_270;
	 wire execution_unit_0_register_file_0_n_178;
	 wire execution_unit_0_register_file_0_n_181;
	 wire execution_unit_0_register_file_0_n_196;
	 wire execution_unit_0_register_file_0_n_179;
	 wire execution_unit_0_register_file_0_n_159;
	 wire execution_unit_0_register_file_0_n_162;
	 wire execution_unit_0_register_file_0_n_177;
	 wire execution_unit_0_register_file_0_n_160;
	 wire execution_unit_0_register_file_0_n_140;
	 wire execution_unit_0_register_file_0_n_143;
	 wire execution_unit_0_register_file_0_n_158;
	 wire execution_unit_0_register_file_0_n_141;
	 wire execution_unit_0_register_file_0_n_121;
	 wire execution_unit_0_register_file_0_n_124;
	 wire execution_unit_0_register_file_0_n_139;
	 wire execution_unit_0_register_file_0_n_122;
	 wire execution_unit_0_register_file_0_n_102;
	 wire execution_unit_0_register_file_0_n_105;
	 wire execution_unit_0_register_file_0_n_120;
	 wire execution_unit_0_register_file_0_n_103;
	 wire execution_unit_0_register_file_0_n_83;
	 wire execution_unit_0_register_file_0_n_86;
	 wire execution_unit_0_register_file_0_n_101;
	 wire execution_unit_0_register_file_0_n_84;
	 wire execution_unit_0_register_file_0_n_64;
	 wire execution_unit_0_register_file_0_n_67;
	 wire execution_unit_0_register_file_0_n_82;
	 wire execution_unit_0_register_file_0_n_65;
	 wire execution_unit_0_register_file_0_n_45;
	 wire execution_unit_0_register_file_0_n_48;
	 wire execution_unit_0_register_file_0_n_63;
	 wire execution_unit_0_register_file_0_n_46;
	 wire execution_unit_0_register_file_0_n_197;
	 wire execution_unit_0_register_file_0_n_200;
	 wire execution_unit_0_register_file_0_n_215;
	 wire execution_unit_0_register_file_0_n_198;
	 wire execution_unit_0_register_file_0_n_254;
	 wire execution_unit_0_register_file_0_n_235;
	 wire execution_unit_0_register_file_0_n_238;
	 wire execution_unit_0_register_file_0_n_253;
	 wire execution_unit_0_register_file_0_n_236;
	 wire execution_unit_0_register_file_0_n_216;
	 wire execution_unit_0_register_file_0_n_219;
	 wire execution_unit_0_register_file_0_n_234;
	 wire execution_unit_0_register_file_0_n_217;
	 wire execution_unit_0_register_file_0_n_28;
	 wire execution_unit_0_register_file_0_n_9;
	 wire execution_unit_0_register_file_0_n_13;
	 wire execution_unit_0_register_file_0_n_180;
	 wire execution_unit_0_register_file_0_n_161;
	 wire execution_unit_0_register_file_0_n_142;
	 wire execution_unit_0_register_file_0_n_123;
	 wire execution_unit_0_register_file_0_n_104;
	 wire execution_unit_0_register_file_0_n_85;
	 wire execution_unit_0_register_file_0_n_66;
	 wire execution_unit_0_register_file_0_n_47;
	 wire execution_unit_0_register_file_0_n_199;
	 wire execution_unit_0_register_file_0_n_237;
	 wire execution_unit_0_register_file_0_n_218;
	 wire execution_unit_0_register_file_0_n_30;
	 wire execution_unit_0_register_file_0_n_11;
	 wire execution_unit_0_register_file_0_n_15;
	 wire execution_unit_0_register_file_0_n_256;
	 wire execution_unit_0_register_file_0_n_274;
	 wire execution_unit_0_register_file_0_n_182;
	 wire execution_unit_0_register_file_0_n_163;
	 wire execution_unit_0_register_file_0_n_144;
	 wire execution_unit_0_register_file_0_n_125;
	 wire execution_unit_0_register_file_0_n_106;
	 wire execution_unit_0_register_file_0_n_87;
	 wire execution_unit_0_register_file_0_n_68;
	 wire execution_unit_0_register_file_0_n_49;
	 wire execution_unit_0_register_file_0_n_201;
	 wire execution_unit_0_register_file_0_n_239;
	 wire execution_unit_0_register_file_0_n_220;
	 wire execution_unit_0_register_file_0_n_257;
	 wire execution_unit_0_register_file_0_n_275;
	 wire execution_unit_0_register_file_0_n_183;
	 wire execution_unit_0_register_file_0_n_164;
	 wire execution_unit_0_register_file_0_n_145;
	 wire execution_unit_0_register_file_0_n_126;
	 wire execution_unit_0_register_file_0_n_107;
	 wire execution_unit_0_register_file_0_n_88;
	 wire execution_unit_0_register_file_0_n_69;
	 wire execution_unit_0_register_file_0_n_50;
	 wire execution_unit_0_register_file_0_n_202;
	 wire execution_unit_0_register_file_0_n_240;
	 wire execution_unit_0_register_file_0_n_221;
	 wire execution_unit_0_register_file_0_n_32;
	 wire execution_unit_0_register_file_0_n_258;
	 wire execution_unit_0_register_file_0_n_276;
	 wire execution_unit_0_register_file_0_n_184;
	 wire execution_unit_0_register_file_0_n_165;
	 wire execution_unit_0_register_file_0_n_146;
	 wire execution_unit_0_register_file_0_n_127;
	 wire execution_unit_0_register_file_0_n_108;
	 wire execution_unit_0_register_file_0_n_89;
	 wire execution_unit_0_register_file_0_n_70;
	 wire execution_unit_0_register_file_0_n_51;
	 wire execution_unit_0_register_file_0_n_203;
	 wire execution_unit_0_register_file_0_n_241;
	 wire execution_unit_0_register_file_0_n_222;
	 wire execution_unit_0_register_file_0_n_259;
	 wire execution_unit_0_register_file_0_n_277;
	 wire execution_unit_0_register_file_0_n_185;
	 wire execution_unit_0_register_file_0_n_166;
	 wire execution_unit_0_register_file_0_n_147;
	 wire execution_unit_0_register_file_0_n_128;
	 wire execution_unit_0_register_file_0_n_109;
	 wire execution_unit_0_register_file_0_n_90;
	 wire execution_unit_0_register_file_0_n_71;
	 wire execution_unit_0_register_file_0_n_52;
	 wire execution_unit_0_register_file_0_n_204;
	 wire execution_unit_0_register_file_0_n_242;
	 wire execution_unit_0_register_file_0_n_223;
	 wire execution_unit_0_register_file_0_n_34;
	 wire execution_unit_0_register_file_0_n_18;
	 wire execution_unit_0_register_file_0_n_260;
	 wire execution_unit_0_register_file_0_n_278;
	 wire execution_unit_0_register_file_0_n_186;
	 wire execution_unit_0_register_file_0_n_167;
	 wire execution_unit_0_register_file_0_n_148;
	 wire execution_unit_0_register_file_0_n_129;
	 wire execution_unit_0_register_file_0_n_110;
	 wire execution_unit_0_register_file_0_n_91;
	 wire execution_unit_0_register_file_0_n_72;
	 wire execution_unit_0_register_file_0_n_53;
	 wire execution_unit_0_register_file_0_n_205;
	 wire execution_unit_0_register_file_0_n_243;
	 wire execution_unit_0_register_file_0_n_224;
	 wire execution_unit_0_register_file_0_n_261;
	 wire execution_unit_0_register_file_0_n_279;
	 wire execution_unit_0_register_file_0_n_187;
	 wire execution_unit_0_register_file_0_n_168;
	 wire execution_unit_0_register_file_0_n_149;
	 wire execution_unit_0_register_file_0_n_130;
	 wire execution_unit_0_register_file_0_n_111;
	 wire execution_unit_0_register_file_0_n_92;
	 wire execution_unit_0_register_file_0_n_73;
	 wire execution_unit_0_register_file_0_n_54;
	 wire execution_unit_0_register_file_0_n_206;
	 wire execution_unit_0_register_file_0_n_244;
	 wire execution_unit_0_register_file_0_n_225;
	 wire execution_unit_0_register_file_0_n_36;
	 wire execution_unit_0_register_file_0_n_12;
	 wire execution_unit_0_register_file_0_n_20;
	 wire execution_unit_0_register_file_0_n_262;
	 wire execution_unit_0_register_file_0_n_280;
	 wire execution_unit_0_register_file_0_n_188;
	 wire execution_unit_0_register_file_0_n_169;
	 wire execution_unit_0_register_file_0_n_150;
	 wire execution_unit_0_register_file_0_n_131;
	 wire execution_unit_0_register_file_0_n_112;
	 wire execution_unit_0_register_file_0_n_93;
	 wire execution_unit_0_register_file_0_n_74;
	 wire execution_unit_0_register_file_0_n_55;
	 wire execution_unit_0_register_file_0_n_207;
	 wire execution_unit_0_register_file_0_n_245;
	 wire execution_unit_0_register_file_0_n_226;
	 wire execution_unit_0_register_file_0_n_263;
	 wire execution_unit_0_register_file_0_n_281;
	 wire execution_unit_0_register_file_0_n_189;
	 wire execution_unit_0_register_file_0_n_170;
	 wire execution_unit_0_register_file_0_n_151;
	 wire execution_unit_0_register_file_0_n_132;
	 wire execution_unit_0_register_file_0_n_113;
	 wire execution_unit_0_register_file_0_n_94;
	 wire execution_unit_0_register_file_0_n_75;
	 wire execution_unit_0_register_file_0_n_56;
	 wire execution_unit_0_register_file_0_n_208;
	 wire execution_unit_0_register_file_0_n_246;
	 wire execution_unit_0_register_file_0_n_227;
	 wire execution_unit_0_register_file_0_n_38;
	 wire execution_unit_0_register_file_0_n_5;
	 wire execution_unit_0_register_file_0_n_264;
	 wire execution_unit_0_register_file_0_n_282;
	 wire execution_unit_0_register_file_0_n_190;
	 wire execution_unit_0_register_file_0_n_171;
	 wire execution_unit_0_register_file_0_n_152;
	 wire execution_unit_0_register_file_0_n_133;
	 wire execution_unit_0_register_file_0_n_114;
	 wire execution_unit_0_register_file_0_n_95;
	 wire execution_unit_0_register_file_0_n_76;
	 wire execution_unit_0_register_file_0_n_57;
	 wire execution_unit_0_register_file_0_n_209;
	 wire execution_unit_0_register_file_0_n_247;
	 wire execution_unit_0_register_file_0_n_228;
	 wire execution_unit_0_register_file_0_n_265;
	 wire execution_unit_0_register_file_0_n_283;
	 wire execution_unit_0_register_file_0_n_191;
	 wire execution_unit_0_register_file_0_n_172;
	 wire execution_unit_0_register_file_0_n_153;
	 wire execution_unit_0_register_file_0_n_134;
	 wire execution_unit_0_register_file_0_n_115;
	 wire execution_unit_0_register_file_0_n_96;
	 wire execution_unit_0_register_file_0_n_77;
	 wire execution_unit_0_register_file_0_n_58;
	 wire execution_unit_0_register_file_0_n_210;
	 wire execution_unit_0_register_file_0_n_248;
	 wire execution_unit_0_register_file_0_n_229;
	 wire execution_unit_0_register_file_0_n_40;
	 wire execution_unit_0_register_file_0_n_3;
	 wire execution_unit_0_register_file_0_n_266;
	 wire execution_unit_0_register_file_0_n_284;
	 wire execution_unit_0_register_file_0_n_192;
	 wire execution_unit_0_register_file_0_n_173;
	 wire execution_unit_0_register_file_0_n_154;
	 wire execution_unit_0_register_file_0_n_135;
	 wire execution_unit_0_register_file_0_n_116;
	 wire execution_unit_0_register_file_0_n_97;
	 wire execution_unit_0_register_file_0_n_78;
	 wire execution_unit_0_register_file_0_n_59;
	 wire execution_unit_0_register_file_0_n_211;
	 wire execution_unit_0_register_file_0_n_249;
	 wire execution_unit_0_register_file_0_n_230;
	 wire execution_unit_0_register_file_0_n_267;
	 wire execution_unit_0_register_file_0_n_285;
	 wire execution_unit_0_register_file_0_n_193;
	 wire execution_unit_0_register_file_0_n_174;
	 wire execution_unit_0_register_file_0_n_155;
	 wire execution_unit_0_register_file_0_n_136;
	 wire execution_unit_0_register_file_0_n_117;
	 wire execution_unit_0_register_file_0_n_98;
	 wire execution_unit_0_register_file_0_n_79;
	 wire execution_unit_0_register_file_0_n_60;
	 wire execution_unit_0_register_file_0_n_212;
	 wire execution_unit_0_register_file_0_n_250;
	 wire execution_unit_0_register_file_0_n_231;
	 wire execution_unit_0_register_file_0_n_42;
	 wire execution_unit_0_register_file_0_n_1;
	 wire execution_unit_0_register_file_0_n_268;
	 wire execution_unit_0_register_file_0_n_286;
	 wire execution_unit_0_register_file_0_n_194;
	 wire execution_unit_0_register_file_0_n_175;
	 wire execution_unit_0_register_file_0_n_156;
	 wire execution_unit_0_register_file_0_n_137;
	 wire execution_unit_0_register_file_0_n_118;
	 wire execution_unit_0_register_file_0_n_99;
	 wire execution_unit_0_register_file_0_n_80;
	 wire execution_unit_0_register_file_0_n_61;
	 wire execution_unit_0_register_file_0_n_213;
	 wire execution_unit_0_register_file_0_n_251;
	 wire execution_unit_0_register_file_0_n_232;
	 wire execution_unit_0_register_file_0_n_269;
	 wire execution_unit_0_register_file_0_n_287;
	 wire execution_unit_0_register_file_0_n_195;
	 wire execution_unit_0_register_file_0_n_176;
	 wire execution_unit_0_register_file_0_n_157;
	 wire execution_unit_0_register_file_0_n_138;
	 wire execution_unit_0_register_file_0_n_119;
	 wire execution_unit_0_register_file_0_n_100;
	 wire execution_unit_0_register_file_0_n_81;
	 wire execution_unit_0_register_file_0_n_62;
	 wire execution_unit_0_register_file_0_n_214;
	 wire execution_unit_0_register_file_0_n_252;
	 wire execution_unit_0_register_file_0_n_233;
	 wire execution_unit_0_register_file_0_n_43;
	 wire clock_module_0_cpuoff_and_mclk_dma_wkup;
	 wire clock_module_0_cpuoff_and_mclk_dma_wkup_s;
	 wire clock_module_0_mclk_wkup_s;
	 wire clock_module_0_cpuoff_and_mclk_dma_enable;
	 wire clock_module_0_por_noscan;
	 wire clock_module_0_puc_a_scan;
	 wire clock_module_0_puc_noscan_n;
	 wire clock_module_0_scg0_and_mclk_dma_enable;
	 wire clock_module_0_cpuoff_and_mclk_enable;
	 wire clock_module_0_cpu_enabled_with_dco;
	 wire clock_module_0_dco_not_enabled_by_dbg;
	 wire clock_module_0_dco_disable_by_scg0;
	 wire clock_module_0_dco_disable_by_cpu_en;
	 wire clock_module_0_dco_enable_nxt;
	 wire clock_module_0_scg0_and_mclk_dma_wkup;
	 wire clock_module_0_dco_en_wkup;
	 wire clock_module_0_dco_mclk_wkup;
	 wire clock_module_0_dco_wkup_set_scan_observe;
	 wire clock_module_0_dco_wkup_set_scan;
	 wire clock_module_0_dco_wkup_n;
	 wire clock_module_0_scg1_and_mclk_dma_enable;
	 wire clock_module_0_scg1_and_mclk_dma_wkup;
	 wire clock_module_0_scg1_and_mclk_dma_wkup_s;
	 wire clock_module_0_nodiv_mclk_n;
	 wire clock_module_0_dco_disable;
	 wire clock_module_0_n_1_0;
	 wire clock_module_0_n_7_0;
	 wire clock_module_0_n_7_1;
	 wire clock_module_0_n_7_2;
	 wire clock_module_0_n_7_3;
	 wire clock_module_0_reg_sel;
	 wire clock_module_0_reg_read;
	 wire clock_module_0_n_10_0;
	 wire clock_module_0_n_11_0;
	 wire clock_module_0_reg_lo_write;
	 wire clock_module_0_bcsctl2_wr;
	 wire [7:0]clock_module_0_bcsctl2;
	 wire clock_module_0_reg_hi_write;
	 wire clock_module_0_bcsctl1_wr;
	 wire [7:0]clock_module_0_bcsctl1;
	 wire [2:0]clock_module_0_aclk_div;
	 wire clock_module_0_n_23_0;
	 wire clock_module_0_n_23_1;
	 wire clock_module_0_n_28_0;
	 wire clock_module_0_n_28_1;
	 wire clock_module_0_n_28_2;
	 wire clock_module_0_n_28_3;
	 wire clock_module_0_n_28_4;
	 wire clock_module_0_n_28_5;
	 wire clock_module_0_n_28_6;
	 wire clock_module_0_n_28_7;
	 wire clock_module_0_n_28_8;
	 wire clock_module_0_n_28_9;
	 wire clock_module_0_aclk_div_sel;
	 wire clock_module_0_n_29_0;
	 wire clock_module_0_aclk_div_en;
	 wire [2:0]clock_module_0_mclk_div;
	 wire clock_module_0_n_31_0;
	 wire clock_module_0_n_31_1;
	 wire clock_module_0_n_36_0;
	 wire clock_module_0_n_36_1;
	 wire clock_module_0_n_36_2;
	 wire clock_module_0_n_36_3;
	 wire clock_module_0_n_36_4;
	 wire clock_module_0_n_36_5;
	 wire clock_module_0_n_36_6;
	 wire clock_module_0_n_36_7;
	 wire clock_module_0_n_36_8;
	 wire clock_module_0_n_36_9;
	 wire clock_module_0_mclk_div_sel;
	 wire clock_module_0_n_37_0;
	 wire clock_module_0_n_37_1;
	 wire clock_module_0_mclk_active;
	 wire clock_module_0_mclk_div_en;
	 wire clock_module_0_n_39_0;
	 wire clock_module_0_mclk_dma_div_en;
	 wire clock_module_0_por_a;
	 wire clock_module_0_dbg_rst_nxt;
	 wire clock_module_0_dbg_rst_noscan;
	 wire clock_module_0_dco_wkup_set;
	 wire clock_module_0_n_46_0;
	 wire [2:0]clock_module_0_smclk_div;
	 wire clock_module_0_n_48_0;
	 wire clock_module_0_n_48_1;
	 wire clock_module_0_n_53_0;
	 wire clock_module_0_n_53_1;
	 wire clock_module_0_n_53_2;
	 wire clock_module_0_n_53_3;
	 wire clock_module_0_n_53_4;
	 wire clock_module_0_n_53_5;
	 wire clock_module_0_n_53_6;
	 wire clock_module_0_n_53_7;
	 wire clock_module_0_n_53_8;
	 wire clock_module_0_n_53_9;
	 wire clock_module_0_smclk_div_sel;
	 wire clock_module_0_n_54_0;
	 wire clock_module_0_n_54_1;
	 wire clock_module_0_n_54_2;
	 wire clock_module_0_smclk_div_en;
	 wire clock_module_0_puc_a;
	 wire clock_module_0_n_5;
	 wire clock_module_0_n_4;
	 wire clock_module_0_n_8;
	 wire clock_module_0_n_10;
	 wire clock_module_0_n_19;
	 wire clock_module_0_n_22;
	 wire clock_module_0_n_18;
	 wire clock_module_0_n_20;
	 wire clock_module_0_n_21;
	 wire clock_module_0_n_23;
	 wire clock_module_0_n_24;
	 wire clock_module_0_n_1;
	 wire clock_module_0_n_28;
	 wire clock_module_0_n_9;
	 wire clock_module_0_n_12;
	 wire clock_module_0_n_15;
	 wire clock_module_0_n_11;
	 wire clock_module_0_n_13;
	 wire clock_module_0_n_14;
	 wire clock_module_0_n_16;
	 wire clock_module_0_n_17;
	 wire clock_module_0_n_39;
	 wire clock_module_0_n_38;
	 wire clock_module_0_n_40;
	 wire clock_module_0_n_25;
	 wire clock_module_0_n_36;
	 wire clock_module_0_n_37;
	 wire clock_module_0_n_26;
	 wire clock_module_0_n_0;
	 wire clock_module_0_n_2;
	 wire clock_module_0_n_41;
	 wire clock_module_0_n_27;
	 wire clock_module_0_n_3;
	 wire clock_module_0_n_6;
	 wire clock_module_0_n_7;
	 wire clock_module_0_n_30;
	 wire clock_module_0_n_33;
	 wire clock_module_0_n_29;
	 wire clock_module_0_n_31;
	 wire clock_module_0_n_32;
	 wire clock_module_0_n_34;
	 wire clock_module_0_n_35;
	 wire clock_module_0_sync_cell_mclk_wkup_n_0;
	 wire clock_module_0_sync_cell_mclk_wkup_n_1;
	 wire clock_module_0_clock_gate_mclk_enable_in;
	 wire clock_module_0_clock_gate_mclk_enable_latch;
	 wire clock_module_0_clock_gate_mclk_n_0;
	 wire clock_module_0_sync_reset_por_n_0;
	 wire clock_module_0_sync_reset_por_n_1;
	 wire clock_module_0_scan_mux_por_n_0_0;
	 wire clock_module_0_scan_mux_por_n_0_1;
	 wire clock_module_0_scan_mux_puc_rst_a_n_0_0;
	 wire clock_module_0_scan_mux_puc_rst_a_n_0_1;
	 wire clock_module_0_sync_cell_puc_n_0;
	 wire clock_module_0_sync_cell_puc_n_1;
	 wire clock_module_0_scan_mux_puc_rst_n_0_0;
	 wire clock_module_0_scan_mux_puc_rst_n_0_1;
	 wire clock_module_0_sync_cell_mclk_dma_wkup_n_0;
	 wire clock_module_0_sync_cell_mclk_dma_wkup_n_1;
	 wire clock_module_0_clock_gate_dma_mclk_enable_in;
	 wire clock_module_0_clock_gate_dma_mclk_enable_latch;
	 wire clock_module_0_clock_gate_dma_mclk_n_0;
	 wire clock_module_0_clock_gate_aclk_enable_in;
	 wire clock_module_0_clock_gate_aclk_enable_latch;
	 wire clock_module_0_clock_gate_aclk_n_0;
	 wire clock_module_0_clock_gate_dbg_clk_enable_in;
	 wire clock_module_0_clock_gate_dbg_clk_enable_latch;
	 wire clock_module_0_clock_gate_dbg_clk_n_0;
	 wire clock_module_0_scan_mux_dbg_rst_n_0_0;
	 wire clock_module_0_scan_mux_dbg_rst_n_0_1;
	 wire clock_module_0_scan_mux_dco_wkup_observe_n_0_0;
	 wire clock_module_0_scan_mux_dco_wkup_observe_n_0_1;
	 wire clock_module_0_scan_mux_dco_wkup_n_0_0;
	 wire clock_module_0_scan_mux_dco_wkup_n_0_1;
	 wire clock_module_0_sync_cell_dco_wkup_n_0;
	 wire clock_module_0_sync_cell_dco_wkup_n_1;
	 wire clock_module_0_sync_cell_smclk_dma_wkup_n_0;
	 wire clock_module_0_sync_cell_smclk_dma_wkup_n_1;
	 wire clock_module_0_clock_gate_smclk_enable_in;
	 wire clock_module_0_clock_gate_smclk_enable_latch;
	 wire clock_module_0_clock_gate_smclk_n_0;


	NOR2_X1_LVT watchdog_0i_1_0 (.A1(per_we[0]),.A2(per_we[1]),.ZN(watchdog_0_n_1));
	NAND3_X1_LVT watchdog_0i_0_0 (.A1(per_addr[4]),.A2(per_addr[7]),.A3(per_en),.ZN(watchdog_0_n_0_0));
	NOR4_X1_LVT watchdog_0i_0_1 (.A1(watchdog_0_n_0_0),.A2(per_addr[12]),.A3(per_addr[13]),.A4(per_addr[0]),.ZN(watchdog_0_n_0_1));
	NOR4_X1_LVT watchdog_0i_0_2 (.A1(per_addr[2]),.A2(per_addr[3]),.A3(per_addr[5]),.A4(per_addr[6]),.ZN(watchdog_0_n_0_2));
	NOR4_X1_LVT watchdog_0i_0_3 (.A1(per_addr[8]),.A2(per_addr[9]),.A3(per_addr[10]),.A4(per_addr[11]),.ZN(watchdog_0_n_0_3));
	NAND3_X1_LVT watchdog_0i_0_4 (.A1(watchdog_0_n_0_1),.A2(watchdog_0_n_0_2),.A3(watchdog_0_n_0_3),.ZN(watchdog_0_n_0_4));
	NOR2_X1_LVT watchdog_0i_0_5 (.A1(watchdog_0_n_0_4),.A2(per_addr[1]),.ZN(watchdog_0_n_0));
	AND2_X1_LVT watchdog_0i_2_0 (.A1(watchdog_0_n_1),.A2(watchdog_0_n_0),.ZN(per_dout_wdog[5]));
	OR2_X1_LVT watchdog_0i_3_0 (.A1(per_we[0]),.A2(per_we[1]),.ZN(watchdog_0_n_2));
	AND2_X1_LVT watchdog_0i_4_0 (.A1(watchdog_0_n_2),.A2(watchdog_0_n_0),.ZN(watchdog_0_reg_wr));
	CLKGATETST_X1_LVT watchdog_0clk_gate_wdtctl_reg (.CK(mclk),.E(watchdog_0_reg_wr),.SE(1'b0),.GCK(watchdog_0_n_3));
	INV_X1_LVT watchdog_0i_5_0 (.A(puc_rst),.ZN(watchdog_0_n_4));
	DFFR_X1_LVT watchdog_0wdtctl_reg___05F05b7___05F05d (.D(per_din[7]),.RN(watchdog_0_n_4),.CK(watchdog_0_n_3),.Q(watchdog_0_wdtctl[7]),.QN());
	AND2_X1_LVT watchdog_0i_7_6 (.A1(per_dout_wdog[5]),.A2(watchdog_0_wdtctl[7]),.ZN(per_dout_wdog[7]));
	DFFR_X1_LVT watchdog_0wdtctl_reg___05F05b6___05F05d (.D(per_din[6]),.RN(watchdog_0_n_4),.CK(watchdog_0_n_3),.Q(wdtnmies),.QN());
	AND2_X1_LVT watchdog_0i_7_5 (.A1(per_dout_wdog[5]),.A2(wdtnmies),.ZN(per_dout_wdog[6]));
	DFFR_X1_LVT watchdog_0wdtctl_reg___05F05b4___05F05d (.D(per_din[4]),.RN(watchdog_0_n_4),.CK(watchdog_0_n_3),.Q(watchdog_0_wdtctl[4]),.QN());
	AND2_X1_LVT watchdog_0i_7_4 (.A1(per_dout_wdog[5]),.A2(watchdog_0_wdtctl[4]),.ZN(per_dout_wdog[4]));
	DFFR_X1_LVT watchdog_0wdtctl_reg___05F05b3___05F05d (.D(1'b0),.RN(watchdog_0_n_4),.CK(watchdog_0_n_3),.Q(watchdog_0_wdtctl[3]),.QN());
	AND2_X1_LVT watchdog_0i_7_3 (.A1(per_dout_wdog[5]),.A2(watchdog_0_wdtctl[3]),.ZN(per_dout_wdog[3]));
	DFFR_X1_LVT watchdog_0wdtctl_reg___05F05b2___05F05d (.D(1'b0),.RN(watchdog_0_n_4),.CK(watchdog_0_n_3),.Q(watchdog_0_wdtctl[2]),.QN());
	AND2_X1_LVT watchdog_0i_7_2 (.A1(per_dout_wdog[5]),.A2(watchdog_0_wdtctl[2]),.ZN(per_dout_wdog[2]));
	DFFR_X1_LVT watchdog_0wdtctl_reg___05F05b1___05F05d (.D(per_din[1]),.RN(watchdog_0_n_4),.CK(watchdog_0_n_3),.Q(watchdog_0_wdtctl[1]),.QN());
	AND2_X1_LVT watchdog_0i_7_1 (.A1(per_dout_wdog[5]),.A2(watchdog_0_wdtctl[1]),.ZN(per_dout_wdog[1]));
	DFFR_X1_LVT watchdog_0wdtctl_reg___05F05b0___05F05d (.D(per_din[0]),.RN(watchdog_0_n_4),.CK(watchdog_0_n_3),.Q(watchdog_0_wdtctl[0]),.QN());
	AND2_X1_LVT watchdog_0i_7_0 (.A1(watchdog_0_wdtctl[0]),.A2(per_dout_wdog[5]),.ZN(per_dout_wdog[0]));
	INV_X1_LVT watchdog_0i_32_0 (.A(watchdog_0_wdt_evt_toggle),.ZN(watchdog_0_n_30));
	INV_X1_LVT watchdog_0sync_reset_pori_0_0 (.A(puc_rst),.ZN(watchdog_0_sync_reset_por_n_0));
	DFFS_X1_LVT watchdog_0sync_reset_pordata_sync_reg___05F05b0___05F05d (.D(1'b0),.SN(watchdog_0_sync_reset_por_n_0),.CK(smclk),.Q(watchdog_0_sync_reset_por_n_1),.QN());
	DFFS_X1_LVT watchdog_0sync_reset_pordata_sync_reg___05F05b1___05F05d (.D(watchdog_0_sync_reset_por_n_1),.SN(watchdog_0_sync_reset_por_n_0),.CK(smclk),.Q(watchdog_0_wdt_rst_noscan),.QN());
	INV_X1_LVT watchdog_0scan_mux_wdt_rsti_0_0 (.A(scan_mode),.ZN(watchdog_0_scan_mux_wdt_rst_n_0_0));
	AOI22_X1_LVT watchdog_0scan_mux_wdt_rsti_0_1 (.A1(watchdog_0_scan_mux_wdt_rst_n_0_0),.A2(watchdog_0_wdt_rst_noscan),.B1(puc_rst),.B2(scan_mode),.ZN(watchdog_0_scan_mux_wdt_rst_n_0_1));
	INV_X1_LVT watchdog_0scan_mux_wdt_rsti_0_2 (.A(watchdog_0_scan_mux_wdt_rst_n_0_1),.ZN(watchdog_0_wdt_rst));
	INV_X1_LVT watchdog_0i_30_0 (.A(watchdog_0_wdt_rst),.ZN(watchdog_0_n_29));
	DFFR_X1_LVT watchdog_0wdtisx_s_reg___05F05b0___05F05d (.D(watchdog_0_wdtctl[0]),.RN(watchdog_0_n_29),.CK(smclk),.Q(watchdog_0_wdtisx_s[0]),.QN());
	DFFR_X1_LVT watchdog_0wdtisx_ss_reg___05F05b0___05F05d (.D(watchdog_0_wdtisx_s[0]),.RN(watchdog_0_n_29),.CK(smclk),.Q(watchdog_0_wdtisx_ss[0]),.QN());
	INV_X1_LVT watchdog_0i_28_0 (.A(watchdog_0_wdtisx_ss[0]),.ZN(watchdog_0_n_28_0));
	DFFR_X1_LVT watchdog_0wdtisx_s_reg___05F05b1___05F05d (.D(watchdog_0_wdtctl[1]),.RN(watchdog_0_n_29),.CK(smclk),.Q(watchdog_0_wdtisx_s[1]),.QN());
	DFFR_X1_LVT watchdog_0wdtisx_ss_reg___05F05b1___05F05d (.D(watchdog_0_wdtisx_s[1]),.RN(watchdog_0_n_29),.CK(smclk),.Q(watchdog_0_wdtisx_ss[1]),.QN());
	AND2_X1_LVT watchdog_0i_28_1 (.A1(watchdog_0_n_28_0),.A2(watchdog_0_wdtisx_ss[1]),.ZN(watchdog_0_n_28_1));
	NOR2_X1_LVT watchdog_0i_28_2 (.A1(watchdog_0_n_28_0),.A2(watchdog_0_wdtisx_ss[1]),.ZN(watchdog_0_n_28_2));
	NOR2_X1_LVT watchdog_0i_28_3 (.A1(watchdog_0_wdtisx_ss[0]),.A2(watchdog_0_wdtisx_ss[1]),.ZN(watchdog_0_n_28_3));
	INV_X1_LVT watchdog_0i_40_0 (.A(watchdog_0_wdtcnt_clr_toggle),.ZN(watchdog_0_n_35));
	AND2_X1_LVT watchdog_0i_38_0 (.A1(per_din[3]),.A2(watchdog_0_reg_wr),.ZN(watchdog_0_wdtcnt_clr_detect));
	CLKGATETST_X1_LVT watchdog_0clk_gate_wdtcnt_clr_toggle_reg (.CK(mclk),.E(watchdog_0_wdtcnt_clr_detect),.SE(1'b0),.GCK(watchdog_0_n_34));
	DFFR_X1_LVT watchdog_0wdtcnt_clr_toggle_reg (.D(watchdog_0_n_35),.RN(watchdog_0_n_4),.CK(watchdog_0_n_34),.Q(watchdog_0_wdtcnt_clr_toggle),.QN());
	INV_X1_LVT watchdog_0sync_cell_wdtcnt_clri_0_0 (.A(watchdog_0_wdt_rst),.ZN(watchdog_0_sync_cell_wdtcnt_clr_n_0));
	DFFR_X1_LVT watchdog_0sync_cell_wdtcnt_clrdata_sync_reg___05F05b0___05F05d (.D(watchdog_0_wdtcnt_clr_toggle),.RN(watchdog_0_sync_cell_wdtcnt_clr_n_0),.CK(smclk),.Q(watchdog_0_sync_cell_wdtcnt_clr_n_1),.QN());
	DFFR_X1_LVT watchdog_0sync_cell_wdtcnt_clrdata_sync_reg___05F05b1___05F05d (.D(watchdog_0_sync_cell_wdtcnt_clr_n_1),.RN(watchdog_0_sync_cell_wdtcnt_clr_n_0),.CK(smclk),.Q(watchdog_0_wdtcnt_clr_sync),.QN());
	DFFR_X1_LVT watchdog_0wdtcnt_clr_sync_dly_reg (.D(watchdog_0_wdtcnt_clr_sync),.RN(watchdog_0_n_29),.CK(smclk),.Q(watchdog_0_wdtcnt_clr_sync_dly),.QN());
	XOR2_X1_LVT watchdog_0i_19_0 (.A(watchdog_0_wdtcnt_clr_sync),.B(watchdog_0_wdtcnt_clr_sync_dly),.Z(watchdog_0_n_19_0));
	OR2_X1_LVT watchdog_0i_19_1 (.A1(watchdog_0_n_19_0),.A2(watchdog_0_wdtqn_edge),.ZN(watchdog_0_wdtcnt_clr));
	INV_X1_LVT watchdog_0i_21_0 (.A(watchdog_0_wdtcnt_clr),.ZN(watchdog_0_n_21_0));
	AND2_X1_LVT watchdog_0i_21_7 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[6]),.ZN(watchdog_0_n_17));
	INV_X1_LVT watchdog_0i_34_0 (.A(watchdog_0_wdtctl[7]),.ZN(watchdog_0_n_31));
	INV_X1_LVT watchdog_0i_37_0 (.A(watchdog_0_n_31),.ZN(watchdog_0_n_37_0));
	NOR2_X1_LVT watchdog_0i_37_1 (.A1(watchdog_0_n_37_0),.A2(dbg_freeze),.ZN(watchdog_0_n_33));
	INV_X1_LVT watchdog_0sync_cell_wdtcnt_incri_0_0 (.A(watchdog_0_wdt_rst),.ZN(watchdog_0_sync_cell_wdtcnt_incr_n_0));
	DFFR_X1_LVT watchdog_0sync_cell_wdtcnt_incrdata_sync_reg___05F05b0___05F05d (.D(watchdog_0_n_33),.RN(watchdog_0_sync_cell_wdtcnt_incr_n_0),.CK(smclk),.Q(watchdog_0_sync_cell_wdtcnt_incr_n_1),.QN());
	DFFR_X1_LVT watchdog_0sync_cell_wdtcnt_incrdata_sync_reg___05F05b1___05F05d (.D(watchdog_0_sync_cell_wdtcnt_incr_n_1),.RN(watchdog_0_sync_cell_wdtcnt_incr_n_0),.CK(smclk),.Q(watchdog_0_wdtcnt_incr),.QN());
	INV_X1_LVT watchdog_0i_22_1 (.A(watchdog_0_wdtcnt_incr),.ZN(watchdog_0_n_22_1));
	INV_X1_LVT watchdog_0i_22_0 (.A(watchdog_0_wdtcnt_clr),.ZN(watchdog_0_n_22_0));
	NAND2_X1_LVT watchdog_0i_22_2 (.A1(watchdog_0_n_22_1),.A2(watchdog_0_n_22_0),.ZN(watchdog_0_n_27));
	CLKGATETST_X1_LVT watchdog_0clk_gate_wdtcnt_reg (.CK(smclk),.E(watchdog_0_n_27),.SE(1'b0),.GCK(watchdog_0_n_10));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b6___05F05d (.D(watchdog_0_n_17),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[6]),.QN());
	AND2_X1_LVT watchdog_0i_21_6 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[5]),.ZN(watchdog_0_n_16));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b5___05F05d (.D(watchdog_0_n_16),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[5]),.QN());
	AND2_X1_LVT watchdog_0i_21_5 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[4]),.ZN(watchdog_0_n_15));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b4___05F05d (.D(watchdog_0_n_15),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[4]),.QN());
	AND2_X1_LVT watchdog_0i_21_4 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[3]),.ZN(watchdog_0_n_14));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b3___05F05d (.D(watchdog_0_n_14),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[3]),.QN());
	AND2_X1_LVT watchdog_0i_21_3 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[2]),.ZN(watchdog_0_n_13));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b2___05F05d (.D(watchdog_0_n_13),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[2]),.QN());
	AND2_X1_LVT watchdog_0i_21_2 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[1]),.ZN(watchdog_0_n_12));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b1___05F05d (.D(watchdog_0_n_12),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[1]),.QN());
	INV_X1_LVT watchdog_0i_24_0 (.A(watchdog_0_wdtcnt[0]),.ZN(watchdog_0_wdtcnt_nxt[0]));
	AND2_X1_LVT watchdog_0i_21_1 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[0]),.ZN(watchdog_0_n_11));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b0___05F05d (.D(watchdog_0_n_11),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[0]),.QN());
	HA_X1_LVT watchdog_0i_24_1 (.A(watchdog_0_wdtcnt[1]),.B(watchdog_0_wdtcnt[0]),.CO(watchdog_0_n_24_0),.S(watchdog_0_wdtcnt_nxt[1]));
	HA_X1_LVT watchdog_0i_24_2 (.A(watchdog_0_wdtcnt[2]),.B(watchdog_0_n_24_0),.CO(watchdog_0_n_24_1),.S(watchdog_0_wdtcnt_nxt[2]));
	HA_X1_LVT watchdog_0i_24_3 (.A(watchdog_0_wdtcnt[3]),.B(watchdog_0_n_24_1),.CO(watchdog_0_n_24_2),.S(watchdog_0_wdtcnt_nxt[3]));
	HA_X1_LVT watchdog_0i_24_4 (.A(watchdog_0_wdtcnt[4]),.B(watchdog_0_n_24_2),.CO(watchdog_0_n_24_3),.S(watchdog_0_wdtcnt_nxt[4]));
	HA_X1_LVT watchdog_0i_24_5 (.A(watchdog_0_wdtcnt[5]),.B(watchdog_0_n_24_3),.CO(watchdog_0_n_24_4),.S(watchdog_0_wdtcnt_nxt[5]));
	HA_X1_LVT watchdog_0i_24_6 (.A(watchdog_0_wdtcnt[6]),.B(watchdog_0_n_24_4),.CO(watchdog_0_n_24_5),.S(watchdog_0_wdtcnt_nxt[6]));
	INV_X1_LVT watchdog_0i_28_4 (.A(watchdog_0_wdtcnt_nxt[6]),.ZN(watchdog_0_n_28_4));
	OR4_X1_LVT watchdog_0i_28_5 (.A1(watchdog_0_n_28_1),.A2(watchdog_0_n_28_2),.A3(watchdog_0_n_28_3),.A4(watchdog_0_n_28_4),.ZN(watchdog_0_n_28_5));
	AND2_X1_LVT watchdog_0i_21_16 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[15]),.ZN(watchdog_0_n_26));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b15___05F05d (.D(watchdog_0_n_26),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[15]),.QN());
	AND2_X1_LVT watchdog_0i_21_15 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[14]),.ZN(watchdog_0_n_25));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b14___05F05d (.D(watchdog_0_n_25),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[14]),.QN());
	AND2_X1_LVT watchdog_0i_21_14 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[13]),.ZN(watchdog_0_n_24));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b13___05F05d (.D(watchdog_0_n_24),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[13]),.QN());
	AND2_X1_LVT watchdog_0i_21_13 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[12]),.ZN(watchdog_0_n_23));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b12___05F05d (.D(watchdog_0_n_23),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[12]),.QN());
	AND2_X1_LVT watchdog_0i_21_12 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[11]),.ZN(watchdog_0_n_22));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b11___05F05d (.D(watchdog_0_n_22),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[11]),.QN());
	AND2_X1_LVT watchdog_0i_21_11 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[10]),.ZN(watchdog_0_n_21));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b10___05F05d (.D(watchdog_0_n_21),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[10]),.QN());
	AND2_X1_LVT watchdog_0i_21_10 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[9]),.ZN(watchdog_0_n_20));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b9___05F05d (.D(watchdog_0_n_20),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[9]),.QN());
	AND2_X1_LVT watchdog_0i_21_9 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[8]),.ZN(watchdog_0_n_19));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b8___05F05d (.D(watchdog_0_n_19),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[8]),.QN());
	AND2_X1_LVT watchdog_0i_21_8 (.A1(watchdog_0_n_21_0),.A2(watchdog_0_wdtcnt_nxt[7]),.ZN(watchdog_0_n_18));
	DFFR_X1_LVT watchdog_0wdtcnt_reg___05F05b7___05F05d (.D(watchdog_0_n_18),.RN(watchdog_0_n_29),.CK(watchdog_0_n_10),.Q(watchdog_0_wdtcnt[7]),.QN());
	HA_X1_LVT watchdog_0i_24_7 (.A(watchdog_0_wdtcnt[7]),.B(watchdog_0_n_24_5),.CO(watchdog_0_n_24_6),.S(watchdog_0_wdtcnt_nxt[7]));
	HA_X1_LVT watchdog_0i_24_8 (.A(watchdog_0_wdtcnt[8]),.B(watchdog_0_n_24_6),.CO(watchdog_0_n_24_7),.S(watchdog_0_wdtcnt_nxt[8]));
	HA_X1_LVT watchdog_0i_24_9 (.A(watchdog_0_wdtcnt[9]),.B(watchdog_0_n_24_7),.CO(watchdog_0_n_24_8),.S(watchdog_0_wdtcnt_nxt[9]));
	HA_X1_LVT watchdog_0i_24_10 (.A(watchdog_0_wdtcnt[10]),.B(watchdog_0_n_24_8),.CO(watchdog_0_n_24_9),.S(watchdog_0_wdtcnt_nxt[10]));
	HA_X1_LVT watchdog_0i_24_11 (.A(watchdog_0_wdtcnt[11]),.B(watchdog_0_n_24_9),.CO(watchdog_0_n_24_10),.S(watchdog_0_wdtcnt_nxt[11]));
	HA_X1_LVT watchdog_0i_24_12 (.A(watchdog_0_wdtcnt[12]),.B(watchdog_0_n_24_10),.CO(watchdog_0_n_24_11),.S(watchdog_0_wdtcnt_nxt[12]));
	HA_X1_LVT watchdog_0i_24_13 (.A(watchdog_0_wdtcnt[13]),.B(watchdog_0_n_24_11),.CO(watchdog_0_n_24_12),.S(watchdog_0_wdtcnt_nxt[13]));
	HA_X1_LVT watchdog_0i_24_14 (.A(watchdog_0_wdtcnt[14]),.B(watchdog_0_n_24_12),.CO(watchdog_0_n_24_13),.S(watchdog_0_wdtcnt_nxt[14]));
	XNOR2_X1_LVT watchdog_0i_24_15 (.A(watchdog_0_wdtcnt[15]),.B(watchdog_0_n_24_13),.ZN(watchdog_0_n_24_14));
	INV_X1_LVT watchdog_0i_24_16 (.A(watchdog_0_n_24_14),.ZN(watchdog_0_wdtcnt_nxt[15]));
	NAND2_X1_LVT watchdog_0i_28_6 (.A1(watchdog_0_n_28_3),.A2(watchdog_0_wdtcnt_nxt[15]),.ZN(watchdog_0_n_28_6));
	NAND2_X1_LVT watchdog_0i_28_7 (.A1(watchdog_0_n_28_2),.A2(watchdog_0_wdtcnt_nxt[13]),.ZN(watchdog_0_n_28_7));
	NAND2_X1_LVT watchdog_0i_28_8 (.A1(watchdog_0_n_28_1),.A2(watchdog_0_wdtcnt_nxt[9]),.ZN(watchdog_0_n_28_8));
	NAND4_X1_LVT watchdog_0i_28_9 (.A1(watchdog_0_n_28_5),.A2(watchdog_0_n_28_6),.A3(watchdog_0_n_28_7),.A4(watchdog_0_n_28_8),.ZN(watchdog_0_wdtqn_reg));
	AND2_X1_LVT watchdog_0i_29_0 (.A1(watchdog_0_wdtqn_reg),.A2(watchdog_0_wdtcnt_incr),.ZN(watchdog_0_wdtqn_edge));
	CLKGATETST_X1_LVT watchdog_0clk_gate_wdt_evt_toggle_reg (.CK(smclk),.E(watchdog_0_wdtqn_edge),.SE(1'b0),.GCK(watchdog_0_n_28));
	DFFR_X1_LVT watchdog_0wdt_evt_toggle_reg (.D(watchdog_0_n_30),.RN(watchdog_0_n_29),.CK(watchdog_0_n_28),.Q(watchdog_0_wdt_evt_toggle),.QN());
	INV_X1_LVT watchdog_0sync_cell_wdt_evti_0_0 (.A(puc_rst),.ZN(watchdog_0_sync_cell_wdt_evt_n_0));
	DFFR_X1_LVT watchdog_0sync_cell_wdt_evtdata_sync_reg___05F05b0___05F05d (.D(watchdog_0_wdt_evt_toggle),.RN(watchdog_0_sync_cell_wdt_evt_n_0),.CK(mclk),.Q(watchdog_0_sync_cell_wdt_evt_n_1),.QN());
	DFFR_X1_LVT watchdog_0sync_cell_wdt_evtdata_sync_reg___05F05b1___05F05d (.D(watchdog_0_sync_cell_wdt_evt_n_1),.RN(watchdog_0_sync_cell_wdt_evt_n_0),.CK(mclk),.Q(watchdog_0_wdt_evt_toggle_sync),.QN());
	DFFR_X1_LVT watchdog_0wdt_evt_toggle_sync_dly_reg (.D(watchdog_0_wdt_evt_toggle_sync),.RN(watchdog_0_n_4),.CK(mclk),.Q(watchdog_0_wdt_evt_toggle_sync_dly),.QN());
	XOR2_X1_LVT watchdog_0i_9_0 (.A(watchdog_0_wdt_evt_toggle_sync_dly),.B(watchdog_0_wdt_evt_toggle_sync),.Z(watchdog_0_n_9_0));
	INV_X1_LVT watchdog_0i_8_0 (.A(watchdog_0_reg_wr),.ZN(watchdog_0_n_8_0));
	AND4_X1_LVT watchdog_0i_8_1 (.A1(per_din[9]),.A2(per_din[11]),.A3(per_din[12]),.A4(per_din[14]),.ZN(watchdog_0_n_8_1));
	NOR4_X1_LVT watchdog_0i_8_2 (.A1(per_din[8]),.A2(per_din[10]),.A3(per_din[13]),.A4(per_din[15]),.ZN(watchdog_0_n_8_2));
	AOI21_X1_LVT watchdog_0i_8_3 (.A(watchdog_0_n_8_0),.B1(watchdog_0_n_8_1),.B2(watchdog_0_n_8_2),.ZN(watchdog_0_wdtpw_error));
	OR3_X1_LVT watchdog_0i_9_1 (.A1(watchdog_0_n_9_0),.A2(wdtifg_sw_set),.A3(watchdog_0_wdtpw_error),.ZN(watchdog_0_wdtifg_set));
	AOI21_X1_LVT watchdog_0i_10_0 (.A(wdtifg_sw_clr),.B1(irq_acc[10]),.B2(watchdog_0_wdtctl[4]),.ZN(watchdog_0_n_10_0));
	INV_X1_LVT watchdog_0i_10_1 (.A(watchdog_0_n_10_0),.ZN(watchdog_0_wdtifg_clr));
	INV_X1_LVT watchdog_0i_13_1 (.A(watchdog_0_wdtifg_clr),.ZN(watchdog_0_n_13_1));
	INV_X1_LVT watchdog_0i_13_0 (.A(watchdog_0_wdtifg_set),.ZN(watchdog_0_n_13_0));
	NAND2_X1_LVT watchdog_0i_13_2 (.A1(watchdog_0_n_13_1),.A2(watchdog_0_n_13_0),.ZN(watchdog_0_n_7));
	CLKGATETST_X1_LVT watchdog_0clk_gate_wdtifg_reg (.CK(mclk),.E(watchdog_0_n_7),.SE(1'b0),.GCK(watchdog_0_n_5));
	INV_X1_LVT watchdog_0i_11_0 (.A(por),.ZN(watchdog_0_n_6));
	DFFR_X1_LVT watchdog_0wdtifg_reg (.D(watchdog_0_wdtifg_set),.RN(watchdog_0_n_6),.CK(watchdog_0_n_5),.Q(wdtifg),.QN());
	AND3_X1_LVT watchdog_0i_15_0 (.A1(watchdog_0_wdtctl[4]),.A2(wdtie),.A3(wdtifg),.ZN(wdt_irq));
	INV_X1_LVT watchdog_0i_16_0 (.A(watchdog_0_wdtctl[4]),.ZN(watchdog_0_n_8));
	AOI21_X1_LVT watchdog_0i_17_0 (.A(watchdog_0_wdtpw_error),.B1(watchdog_0_wdtifg_set),.B2(watchdog_0_n_8),.ZN(watchdog_0_n_17_0));
	INV_X1_LVT watchdog_0i_17_1 (.A(watchdog_0_n_17_0),.ZN(watchdog_0_n_9));
	DFFR_X1_LVT watchdog_0wdt_reset_reg (.D(watchdog_0_n_9),.RN(watchdog_0_n_6),.CK(mclk),.Q(wdt_reset),.QN());
	DFFS_X1_LVT watchdog_0wdtifg_clr_reg_reg (.D(watchdog_0_wdtifg_clr),.SN(watchdog_0_n_4),.CK(mclk),.Q(watchdog_0_wdtifg_clr_reg),.QN());
	DFFR_X1_LVT watchdog_0wdtqn_edge_reg_reg (.D(watchdog_0_wdtqn_edge),.RN(watchdog_0_n_29),.CK(smclk),.Q(watchdog_0_wdtqn_edge_reg),.QN());
	INV_X1_LVT watchdog_0wakeup_cell_wdogscan_mux_clki_0_0 (.A(scan_mode),.ZN(watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_0));
	AOI22_X1_LVT watchdog_0wakeup_cell_wdogscan_mux_clki_0_1 (.A1(watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_0),.A2(watchdog_0_wdtqn_edge_reg),.B1(mclk),.B2(scan_mode),.ZN(watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_1));
	INV_X1_LVT watchdog_0wakeup_cell_wdogscan_mux_clki_0_2 (.A(watchdog_0_wakeup_cell_wdog_scan_mux_clk_n_0_1),.ZN(watchdog_0_wakeup_cell_wdog_wkup_clk));
	INV_X1_LVT watchdog_0wakeup_cell_wdogscan_mux_rsti_0_0 (.A(scan_mode),.ZN(watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_0));
	AOI22_X1_LVT watchdog_0wakeup_cell_wdogscan_mux_rsti_0_1 (.A1(watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_0),.A2(watchdog_0_wdtifg_clr_reg),.B1(puc_rst),.B2(scan_mode),.ZN(watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_1));
	INV_X1_LVT watchdog_0wakeup_cell_wdogscan_mux_rsti_0_2 (.A(watchdog_0_wakeup_cell_wdog_scan_mux_rst_n_0_1),.ZN(watchdog_0_wakeup_cell_wdog_wkup_rst));
	INV_X1_LVT watchdog_0wakeup_cell_wdogi_0_0 (.A(watchdog_0_wakeup_cell_wdog_wkup_rst),.ZN(watchdog_0_wakeup_cell_wdog_n_0));
	DFFR_X1_LVT watchdog_0wakeup_cell_wdogwkup_out_reg (.D(1'b1),.RN(watchdog_0_wakeup_cell_wdog_n_0),.CK(watchdog_0_wakeup_cell_wdog_wkup_clk),.Q(watchdog_0_wdt_wkup_pre),.QN());
	NOR2_X1_LVT watchdog_0i_35_2 (.A1(wdtie),.A2(watchdog_0_n_8),.ZN(watchdog_0_n_35_1));
	INV_X1_LVT watchdog_0i_35_0 (.A(watchdog_0_n_31),.ZN(watchdog_0_n_35_0));
	NOR2_X1_LVT watchdog_0i_35_1 (.A1(watchdog_0_n_35_1),.A2(watchdog_0_n_35_0),.ZN(watchdog_0_n_32));
	DFFR_X1_LVT watchdog_0wdt_wkup_en_reg (.D(watchdog_0_n_32),.RN(watchdog_0_n_4),.CK(mclk),.Q(watchdog_0_wdt_wkup_en),.QN());
	AND2_X1_LVT watchdog_0and_wdt_wkupi_0_0 (.A1(watchdog_0_wdt_wkup_pre),.A2(watchdog_0_wdt_wkup_en),.ZN(wdt_wkup));
	DFFR_X1_LVT watchdog_0wdtctl_reg___05F05b5___05F05d (.D(1'b0),.RN(watchdog_0_n_4),.CK(watchdog_0_n_3),.Q(watchdog_0_wdtctl[5]),.QN());
	INV_X1_LVT sfr_0i_13_1 (.A(per_din[4]),.ZN(sfr_0_n_13_1));
	INV_X1_LVT sfr_0i_0_0 (.A(per_en),.ZN(sfr_0_n_0_0));
	NOR4_X1_LVT sfr_0i_0_1 (.A1(sfr_0_n_0_0),.A2(per_addr[11]),.A3(per_addr[12]),.A4(per_addr[13]),.ZN(sfr_0_n_0_1));
	NOR4_X1_LVT sfr_0i_0_2 (.A1(per_addr[3]),.A2(per_addr[4]),.A3(per_addr[5]),.A4(per_addr[6]),.ZN(sfr_0_n_0_2));
	NOR4_X1_LVT sfr_0i_0_3 (.A1(per_addr[7]),.A2(per_addr[8]),.A3(per_addr[9]),.A4(per_addr[10]),.ZN(sfr_0_n_0_3));
	AND3_X1_LVT sfr_0i_0_4 (.A1(sfr_0_n_0_1),.A2(sfr_0_n_0_2),.A3(sfr_0_n_0_3),.ZN(sfr_0_reg_sel));
	AND2_X1_LVT sfr_0i_1_0 (.A1(per_we[0]),.A2(sfr_0_reg_sel),.ZN(sfr_0_reg_lo_write));
	INV_X1_LVT sfr_0i_2_1 (.A(per_addr[1]),.ZN(sfr_0_n_2_1));
	NAND2_X1_LVT sfr_0i_2_3 (.A1(per_addr[0]),.A2(sfr_0_n_2_1),.ZN(sfr_0_n_2_3));
	NOR2_X1_LVT sfr_0i_2_8 (.A1(sfr_0_n_2_3),.A2(per_addr[2]),.ZN(sfr_0_n_1));
	AND2_X1_LVT sfr_0i_3_1 (.A1(sfr_0_reg_lo_write),.A2(sfr_0_n_1),.ZN(sfr_0_ifg1_wr));
	INV_X1_LVT sfr_0i_4_0 (.A(sfr_0_ifg1_wr),.ZN(sfr_0_n_4_0));
	NOR2_X1_LVT sfr_0i_4_1 (.A1(sfr_0_n_4_0),.A2(per_din[4]),.ZN(sfr_0_n_6));
	INV_X1_LVT sfr_0i_11_0 (.A(puc_rst),.ZN(sfr_0_n_11));
	DFFS_X1_LVT sfr_0nmi_capture_rst_reg (.D(sfr_0_n_6),.SN(sfr_0_n_11),.CK(mclk),.Q(sfr_0_nmi_capture_rst),.QN());
	XOR2_X1_LVT sfr_0i_31_0 (.A(nmi),.B(wdtnmies),.Z(sfr_0_nmi_pol));
	INV_X1_LVT sfr_0wakeup_cell_nmiscan_mux_clki_0_0 (.A(scan_mode),.ZN(sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_0));
	AOI22_X1_LVT sfr_0wakeup_cell_nmiscan_mux_clki_0_1 (.A1(sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_0),.A2(sfr_0_nmi_pol),.B1(mclk),.B2(scan_mode),.ZN(sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_1));
	INV_X1_LVT sfr_0wakeup_cell_nmiscan_mux_clki_0_2 (.A(sfr_0_wakeup_cell_nmi_scan_mux_clk_n_0_1),.ZN(sfr_0_wakeup_cell_nmi_wkup_clk));
	INV_X1_LVT sfr_0wakeup_cell_nmiscan_mux_rsti_0_0 (.A(scan_mode),.ZN(sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_0));
	AOI22_X1_LVT sfr_0wakeup_cell_nmiscan_mux_rsti_0_1 (.A1(sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_0),.A2(sfr_0_nmi_capture_rst),.B1(puc_rst),.B2(scan_mode),.ZN(sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_1));
	INV_X1_LVT sfr_0wakeup_cell_nmiscan_mux_rsti_0_2 (.A(sfr_0_wakeup_cell_nmi_scan_mux_rst_n_0_1),.ZN(sfr_0_wakeup_cell_nmi_wkup_rst));
	INV_X1_LVT sfr_0wakeup_cell_nmii_0_0 (.A(sfr_0_wakeup_cell_nmi_wkup_rst),.ZN(sfr_0_wakeup_cell_nmi_n_0));
	DFFR_X1_LVT sfr_0wakeup_cell_nmiwkup_out_reg (.D(1'b1),.RN(sfr_0_wakeup_cell_nmi_n_0),.CK(sfr_0_wakeup_cell_nmi_wkup_clk),.Q(sfr_0_nmi_capture),.QN());
	INV_X1_LVT sfr_0sync_cell_nmii_0_0 (.A(puc_rst),.ZN(sfr_0_sync_cell_nmi_n_0));
	DFFR_X1_LVT sfr_0sync_cell_nmidata_sync_reg___05F05b0___05F05d (.D(sfr_0_nmi_capture),.RN(sfr_0_sync_cell_nmi_n_0),.CK(mclk),.Q(sfr_0_sync_cell_nmi_n_1),.QN());
	DFFR_X1_LVT sfr_0sync_cell_nmidata_sync_reg___05F05b1___05F05d (.D(sfr_0_sync_cell_nmi_n_1),.RN(sfr_0_sync_cell_nmi_n_0),.CK(mclk),.Q(sfr_0_nmi_s),.QN());
	INV_X1_LVT sfr_0i_10_0 (.A(sfr_0_nmi_s),.ZN(sfr_0_n_10_0));
	DFFR_X1_LVT sfr_0nmi_dly_reg (.D(sfr_0_nmi_s),.RN(sfr_0_n_11),.CK(mclk),.Q(sfr_0_nmi_dly),.QN());
	NOR2_X1_LVT sfr_0i_10_1 (.A1(sfr_0_n_10_0),.A2(sfr_0_nmi_dly),.ZN(sfr_0_nmi_edge));
	INV_X1_LVT sfr_0i_13_0 (.A(sfr_0_nmi_edge),.ZN(sfr_0_n_13_0));
	NAND2_X1_LVT sfr_0i_13_2 (.A1(sfr_0_n_13_1),.A2(sfr_0_n_13_0),.ZN(sfr_0_n_12));
	INV_X1_LVT sfr_0i_14_1 (.A(sfr_0_ifg1_wr),.ZN(sfr_0_n_14_1));
	INV_X1_LVT sfr_0i_14_0 (.A(sfr_0_nmi_edge),.ZN(sfr_0_n_14_0));
	NAND2_X1_LVT sfr_0i_14_2 (.A1(sfr_0_n_14_1),.A2(sfr_0_n_14_0),.ZN(sfr_0_n_13));
	CLKGATETST_X1_LVT sfr_0clk_gate_nmiifg_reg (.CK(mclk),.E(sfr_0_n_13),.SE(1'b0),.GCK(sfr_0_n_10));
	DFFR_X1_LVT sfr_0nmiifg_reg (.D(sfr_0_n_12),.RN(sfr_0_n_11),.CK(sfr_0_n_10),.Q(sfr_0_nmiifg),.QN());
	INV_X1_LVT sfr_0i_7_0 (.A(per_din[4]),.ZN(sfr_0_n_7_0));
	NOR2_X1_LVT sfr_0i_7_1 (.A1(sfr_0_n_7_0),.A2(nmi_acc),.ZN(sfr_0_n_8));
	INV_X1_LVT sfr_0i_2_0 (.A(per_addr[0]),.ZN(sfr_0_n_2_0));
	NAND2_X1_LVT sfr_0i_2_2 (.A1(sfr_0_n_2_0),.A2(sfr_0_n_2_1),.ZN(sfr_0_n_2_2));
	NOR2_X1_LVT sfr_0i_2_7 (.A1(sfr_0_n_2_2),.A2(per_addr[2]),.ZN(sfr_0_n_0));
	AND2_X1_LVT sfr_0i_3_0 (.A1(sfr_0_n_0),.A2(sfr_0_reg_lo_write),.ZN(sfr_0_n_5));
	INV_X1_LVT sfr_0i_8_1 (.A(sfr_0_n_5),.ZN(sfr_0_n_8_1));
	INV_X1_LVT sfr_0i_8_0 (.A(nmi_acc),.ZN(sfr_0_n_8_0));
	NAND2_X1_LVT sfr_0i_8_2 (.A1(sfr_0_n_8_1),.A2(sfr_0_n_8_0),.ZN(sfr_0_n_9));
	CLKGATETST_X1_LVT sfr_0clk_gate_nmie_reg (.CK(mclk),.E(sfr_0_n_9),.SE(1'b0),.GCK(sfr_0_n_7));
	DFFR_X1_LVT sfr_0nmie_reg (.D(sfr_0_n_8),.RN(sfr_0_n_11),.CK(sfr_0_n_7),.Q(sfr_0_nmie),.QN());
	AND2_X1_LVT sfr_0i_16_0 (.A1(sfr_0_nmiifg),.A2(sfr_0_nmie),.ZN(nmi_pnd));
	XOR2_X1_LVT sfr_0i_30_0 (.A(sfr_0_nmi_capture),.B(sfr_0_nmi_dly),.Z(sfr_0_n_31));
	AND2_X1_LVT sfr_0and_nmi_wkupi_0_0 (.A1(sfr_0_n_31),.A2(sfr_0_nmie),.ZN(nmi_wkup));
	NOR2_X1_LVT sfr_0i_17_0 (.A1(per_we[0]),.A2(per_we[1]),.ZN(sfr_0_n_14));
	AND2_X1_LVT sfr_0i_18_0 (.A1(sfr_0_n_14),.A2(sfr_0_reg_sel),.ZN(sfr_0_reg_read));
	INV_X1_LVT sfr_0i_2_6 (.A(per_addr[2]),.ZN(sfr_0_n_2_6));
	NOR2_X1_LVT sfr_0i_2_11 (.A1(sfr_0_n_2_2),.A2(sfr_0_n_2_6),.ZN(sfr_0_n_4));
	AND2_X1_LVT sfr_0i_19_4 (.A1(sfr_0_reg_read),.A2(sfr_0_n_4),.ZN(sfr_0_n_19));
	AND2_X1_LVT sfr_0i_21_7 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(per_dout_sfr[15]));
	AND2_X1_LVT sfr_0i_21_6 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(per_dout_sfr[14]));
	AND2_X1_LVT sfr_0i_21_5 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(per_dout_sfr[13]));
	NAND2_X1_LVT sfr_0i_2_5 (.A1(per_addr[0]),.A2(per_addr[1]),.ZN(sfr_0_n_2_5));
	NOR2_X1_LVT sfr_0i_2_10 (.A1(sfr_0_n_2_5),.A2(per_addr[2]),.ZN(sfr_0_n_3));
	AND2_X1_LVT sfr_0i_19_3 (.A1(sfr_0_reg_read),.A2(sfr_0_n_3),.ZN(sfr_0_n_18));
	AND2_X1_LVT sfr_0i_21_4 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(sfr_0_n_25));
	OR2_X1_LVT sfr_0i_27_6 (.A1(sfr_0_n_18),.A2(sfr_0_n_25),.ZN(per_dout_sfr[12]));
	AND2_X1_LVT sfr_0i_21_3 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(per_dout_sfr[11]));
	AND2_X1_LVT sfr_0i_21_2 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(per_dout_sfr[10]));
	NAND2_X1_LVT sfr_0i_2_4 (.A1(sfr_0_n_2_0),.A2(per_addr[1]),.ZN(sfr_0_n_2_4));
	NOR2_X1_LVT sfr_0i_2_9 (.A1(sfr_0_n_2_4),.A2(per_addr[2]),.ZN(sfr_0_n_2));
	AND2_X1_LVT sfr_0i_19_2 (.A1(sfr_0_reg_read),.A2(sfr_0_n_2),.ZN(sfr_0_n_17));
	AND2_X1_LVT sfr_0i_21_1 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(sfr_0_n_24));
	OR2_X1_LVT sfr_0i_27_5 (.A1(sfr_0_n_17),.A2(sfr_0_n_24),.ZN(per_dout_sfr[9]));
	AND2_X1_LVT sfr_0i_21_0 (.A1(1'b0),.A2(sfr_0_n_19),.ZN(per_dout_sfr[8]));
	AND2_X1_LVT sfr_0i_20_7 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(per_dout_sfr[7]));
	AND2_X1_LVT sfr_0i_20_6 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(per_dout_sfr[6]));
	AND2_X1_LVT sfr_0i_20_5 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(per_dout_sfr[5]));
	AND2_X1_LVT sfr_0i_19_0 (.A1(sfr_0_n_0),.A2(sfr_0_reg_read),.ZN(sfr_0_n_15));
	AND2_X1_LVT sfr_0i_26_0 (.A1(sfr_0_nmie),.A2(sfr_0_n_15),.ZN(sfr_0_n_30));
	AND2_X1_LVT sfr_0i_19_1 (.A1(sfr_0_reg_read),.A2(sfr_0_n_1),.ZN(sfr_0_n_16));
	AND2_X1_LVT sfr_0i_23_0 (.A1(sfr_0_nmiifg),.A2(sfr_0_n_16),.ZN(sfr_0_n_27));
	AND2_X1_LVT sfr_0i_20_4 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(sfr_0_n_23));
	OR4_X1_LVT sfr_0i_27_4 (.A1(sfr_0_n_30),.A2(sfr_0_n_27),.A3(sfr_0_n_18),.A4(sfr_0_n_23),.ZN(per_dout_sfr[4]));
	AND2_X1_LVT sfr_0i_20_3 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(sfr_0_n_22));
	OR2_X1_LVT sfr_0i_27_3 (.A1(sfr_0_n_17),.A2(sfr_0_n_22),.ZN(per_dout_sfr[3]));
	AND2_X1_LVT sfr_0i_20_2 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(per_dout_sfr[2]));
	AND2_X1_LVT sfr_0i_20_1 (.A1(sfr_0_n_19),.A2(1'b0),.ZN(sfr_0_n_21));
	OR2_X1_LVT sfr_0i_27_2 (.A1(sfr_0_n_17),.A2(sfr_0_n_21),.ZN(per_dout_sfr[1]));
	AND2_X1_LVT sfr_0i_22_0 (.A1(wdtifg),.A2(sfr_0_n_16),.ZN(sfr_0_n_26));
	AND2_X1_LVT sfr_0i_20_0 (.A1(1'b0),.A2(sfr_0_n_19),.ZN(sfr_0_n_20));
	OR4_X1_LVT sfr_0i_27_0 (.A1(sfr_0_n_26),.A2(sfr_0_n_17),.A3(sfr_0_n_18),.A4(sfr_0_n_20),.ZN(sfr_0_n_27_0));
	CLKGATETST_X1_LVT sfr_0clk_gate_wdtie_reg (.CK(mclk),.E(sfr_0_n_5),.SE(1'b0),.GCK(sfr_0_n_28));
	DFFR_X1_LVT sfr_0wdtie_reg (.D(per_din[0]),.RN(sfr_0_n_11),.CK(sfr_0_n_28),.Q(wdtie),.QN());
	AND2_X1_LVT sfr_0i_25_0 (.A1(wdtie),.A2(sfr_0_n_15),.ZN(sfr_0_n_29));
	OR2_X1_LVT sfr_0i_27_1 (.A1(sfr_0_n_27_0),.A2(sfr_0_n_29),.ZN(per_dout_sfr[0]));
	INV_X1_LVT sfr_0i_28_0 (.A(sfr_0_ifg1_wr),.ZN(sfr_0_n_28_0));
	NOR2_X1_LVT sfr_0i_28_1 (.A1(sfr_0_n_28_0),.A2(per_din[0]),.ZN(wdtifg_sw_clr));
	AND2_X1_LVT sfr_0i_29_0 (.A1(sfr_0_ifg1_wr),.A2(per_din[0]),.ZN(wdtifg_sw_set));
	INV_X1_LVT dbg_0i_48_2 (.A(dbg_0_dbg_addr[1]),.ZN(dbg_0_n_48_1));
	NAND2_X1_LVT dbg_0i_48_7 (.A1(dbg_0_n_48_1),.A2(dbg_0_n_48_0),.ZN(dbg_0_dbg_addr_in[1]));
	NOR2_X1_LVT dbg_0i_49_2 (.A1(dbg_0_dbg_addr_in[0]),.A2(dbg_0_dbg_addr_in[1]),.ZN(dbg_0_n_49_2));
	INV_X1_LVT dbg_0i_48_3 (.A(dbg_0_dbg_addr[2]),.ZN(dbg_0_n_48_2));
	NAND2_X1_LVT dbg_0i_48_8 (.A1(dbg_0_n_48_2),.A2(dbg_0_n_48_0),.ZN(dbg_0_dbg_addr_in[2]));
	NAND2_X1_LVT dbg_0i_49_11 (.A1(dbg_0_n_49_2),.A2(dbg_0_dbg_addr_in[2]),.ZN(dbg_0_n_49_11));
	AND2_X1_LVT dbg_0i_48_4 (.A1(dbg_0_n_48_0),.A2(dbg_0_dbg_addr[3]),.ZN(dbg_0_dbg_addr_in[3]));
	INV_X1_LVT dbg_0i_49_15 (.A(dbg_0_dbg_addr_in[3]),.ZN(dbg_0_n_49_15));
	AND2_X1_LVT dbg_0i_48_5 (.A1(dbg_0_n_48_0),.A2(dbg_0_dbg_addr[4]),.ZN(dbg_0_dbg_addr_in[4]));
	AND2_X1_LVT dbg_0i_48_6 (.A1(dbg_0_n_48_0),.A2(dbg_0_dbg_addr[5]),.ZN(dbg_0_dbg_addr_in[5]));
	NOR2_X1_LVT dbg_0i_49_16 (.A1(dbg_0_dbg_addr_in[4]),.A2(dbg_0_dbg_addr_in[5]),.ZN(dbg_0_n_49_16));
	NAND2_X1_LVT dbg_0i_49_20 (.A1(dbg_0_n_49_15),.A2(dbg_0_n_49_16),.ZN(dbg_0_n_49_20));
	NOR2_X1_LVT dbg_0i_49_26 (.A1(dbg_0_n_49_11),.A2(dbg_0_n_49_20),.ZN(dbg_0_n_95));
	AND2_X1_LVT dbg_0i_50_2 (.A1(dbg_0_dbg_wr),.A2(dbg_0_n_95),.ZN(dbg_0_mem_ctl_wr));
	AND2_X1_LVT dbg_0i_1_0 (.A1(dbg_0_mem_ctl_wr),.A2(dbg_0_dbg_din[0]),.ZN(dbg_0_n_1));
	INV_X1_LVT dbg_0i_51_0 (.A(dbg_rst),.ZN(dbg_0_n_104));
	DFFR_X1_LVT dbg_0mem_start_reg (.D(dbg_0_n_1),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_start),.QN());
	AND2_X1_LVT dbg_0i_50_5 (.A1(dbg_0_dbg_wr),.A2(dbg_0_n_98),.ZN(dbg_0_n_102));
	INV_X1_LVT dbg_0i_40_0 (.A(dbg_0_n_102),.ZN(dbg_0_n_40_0));
	INV_X1_LVT dbg_0i_39_3 (.A(dbg_0_mem_cnt[0]),.ZN(dbg_0_n_39_2));
	NAND2_X1_LVT dbg_0i_39_2 (.A1(dbg_0_n_55),.A2(dbg_0_n_39_2),.ZN(dbg_0_n_39_1));
	XNOR2_X1_LVT dbg_0i_39_4 (.A(dbg_0_mem_cnt[1]),.B(dbg_0_n_39_1),.ZN(dbg_0_n_57));
	AOI22_X1_LVT dbg_0i_40_3 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_57),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[1]),.ZN(dbg_0_n_40_2));
	INV_X1_LVT dbg_0i_40_4 (.A(dbg_0_n_40_2),.ZN(dbg_0_n_73));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b1___05F05d (.D(dbg_0_n_73),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[1]),.QN());
	OR2_X1_LVT dbg_0i_39_5 (.A1(dbg_0_mem_cnt[1]),.A2(dbg_0_n_39_1),.ZN(dbg_0_n_39_3));
	XNOR2_X1_LVT dbg_0i_39_6 (.A(dbg_0_mem_cnt[2]),.B(dbg_0_n_39_3),.ZN(dbg_0_n_58));
	AOI22_X1_LVT dbg_0i_40_5 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_58),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[2]),.ZN(dbg_0_n_40_3));
	INV_X1_LVT dbg_0i_40_6 (.A(dbg_0_n_40_3),.ZN(dbg_0_n_74));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b2___05F05d (.D(dbg_0_n_74),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[2]),.QN());
	OR2_X1_LVT dbg_0i_39_7 (.A1(dbg_0_mem_cnt[2]),.A2(dbg_0_n_39_3),.ZN(dbg_0_n_39_4));
	XNOR2_X1_LVT dbg_0i_39_8 (.A(dbg_0_mem_cnt[3]),.B(dbg_0_n_39_4),.ZN(dbg_0_n_59));
	AOI22_X1_LVT dbg_0i_40_7 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_59),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[3]),.ZN(dbg_0_n_40_4));
	INV_X1_LVT dbg_0i_40_8 (.A(dbg_0_n_40_4),.ZN(dbg_0_n_75));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b3___05F05d (.D(dbg_0_n_75),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[3]),.QN());
	NOR4_X1_LVT dbg_0i_37_0 (.A1(dbg_0_mem_cnt[0]),.A2(dbg_0_mem_cnt[1]),.A3(dbg_0_mem_cnt[2]),.A4(dbg_0_mem_cnt[3]),.ZN(dbg_0_n_37_0));
	OR2_X1_LVT dbg_0i_39_9 (.A1(dbg_0_mem_cnt[3]),.A2(dbg_0_n_39_4),.ZN(dbg_0_n_39_5));
	XNOR2_X1_LVT dbg_0i_39_10 (.A(dbg_0_mem_cnt[4]),.B(dbg_0_n_39_5),.ZN(dbg_0_n_60));
	AOI22_X1_LVT dbg_0i_40_9 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_60),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[4]),.ZN(dbg_0_n_40_5));
	INV_X1_LVT dbg_0i_40_10 (.A(dbg_0_n_40_5),.ZN(dbg_0_n_76));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b4___05F05d (.D(dbg_0_n_76),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[4]),.QN());
	OR2_X1_LVT dbg_0i_39_11 (.A1(dbg_0_mem_cnt[4]),.A2(dbg_0_n_39_5),.ZN(dbg_0_n_39_6));
	XNOR2_X1_LVT dbg_0i_39_12 (.A(dbg_0_mem_cnt[5]),.B(dbg_0_n_39_6),.ZN(dbg_0_n_61));
	AOI22_X1_LVT dbg_0i_40_11 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_61),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[5]),.ZN(dbg_0_n_40_6));
	INV_X1_LVT dbg_0i_40_12 (.A(dbg_0_n_40_6),.ZN(dbg_0_n_77));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b5___05F05d (.D(dbg_0_n_77),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[5]),.QN());
	OR2_X1_LVT dbg_0i_39_13 (.A1(dbg_0_mem_cnt[5]),.A2(dbg_0_n_39_6),.ZN(dbg_0_n_39_7));
	XNOR2_X1_LVT dbg_0i_39_14 (.A(dbg_0_mem_cnt[6]),.B(dbg_0_n_39_7),.ZN(dbg_0_n_62));
	AOI22_X1_LVT dbg_0i_40_13 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_62),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[6]),.ZN(dbg_0_n_40_7));
	INV_X1_LVT dbg_0i_40_14 (.A(dbg_0_n_40_7),.ZN(dbg_0_n_78));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b6___05F05d (.D(dbg_0_n_78),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[6]),.QN());
	OR2_X1_LVT dbg_0i_39_15 (.A1(dbg_0_mem_cnt[6]),.A2(dbg_0_n_39_7),.ZN(dbg_0_n_39_8));
	XNOR2_X1_LVT dbg_0i_39_16 (.A(dbg_0_mem_cnt[7]),.B(dbg_0_n_39_8),.ZN(dbg_0_n_63));
	AOI22_X1_LVT dbg_0i_40_15 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_63),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[7]),.ZN(dbg_0_n_40_8));
	INV_X1_LVT dbg_0i_40_16 (.A(dbg_0_n_40_8),.ZN(dbg_0_n_79));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b7___05F05d (.D(dbg_0_n_79),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[7]),.QN());
	NOR4_X1_LVT dbg_0i_37_1 (.A1(dbg_0_mem_cnt[4]),.A2(dbg_0_mem_cnt[5]),.A3(dbg_0_mem_cnt[6]),.A4(dbg_0_mem_cnt[7]),.ZN(dbg_0_n_37_1));
	OR2_X1_LVT dbg_0i_39_17 (.A1(dbg_0_mem_cnt[7]),.A2(dbg_0_n_39_8),.ZN(dbg_0_n_39_9));
	XNOR2_X1_LVT dbg_0i_39_18 (.A(dbg_0_mem_cnt[8]),.B(dbg_0_n_39_9),.ZN(dbg_0_n_64));
	AOI22_X1_LVT dbg_0i_40_17 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_64),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[8]),.ZN(dbg_0_n_40_9));
	INV_X1_LVT dbg_0i_40_18 (.A(dbg_0_n_40_9),.ZN(dbg_0_n_80));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b8___05F05d (.D(dbg_0_n_80),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[8]),.QN());
	OR2_X1_LVT dbg_0i_39_19 (.A1(dbg_0_mem_cnt[8]),.A2(dbg_0_n_39_9),.ZN(dbg_0_n_39_10));
	XNOR2_X1_LVT dbg_0i_39_20 (.A(dbg_0_mem_cnt[9]),.B(dbg_0_n_39_10),.ZN(dbg_0_n_65));
	AOI22_X1_LVT dbg_0i_40_19 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_65),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[9]),.ZN(dbg_0_n_40_10));
	INV_X1_LVT dbg_0i_40_20 (.A(dbg_0_n_40_10),.ZN(dbg_0_n_81));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b9___05F05d (.D(dbg_0_n_81),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[9]),.QN());
	OR2_X1_LVT dbg_0i_39_21 (.A1(dbg_0_mem_cnt[9]),.A2(dbg_0_n_39_10),.ZN(dbg_0_n_39_11));
	XNOR2_X1_LVT dbg_0i_39_22 (.A(dbg_0_mem_cnt[10]),.B(dbg_0_n_39_11),.ZN(dbg_0_n_66));
	AOI22_X1_LVT dbg_0i_40_21 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_66),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[10]),.ZN(dbg_0_n_40_11));
	INV_X1_LVT dbg_0i_40_22 (.A(dbg_0_n_40_11),.ZN(dbg_0_n_82));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b10___05F05d (.D(dbg_0_n_82),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[10]),.QN());
	OR2_X1_LVT dbg_0i_39_23 (.A1(dbg_0_mem_cnt[10]),.A2(dbg_0_n_39_11),.ZN(dbg_0_n_39_12));
	XNOR2_X1_LVT dbg_0i_39_24 (.A(dbg_0_mem_cnt[11]),.B(dbg_0_n_39_12),.ZN(dbg_0_n_67));
	AOI22_X1_LVT dbg_0i_40_23 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_67),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[11]),.ZN(dbg_0_n_40_12));
	INV_X1_LVT dbg_0i_40_24 (.A(dbg_0_n_40_12),.ZN(dbg_0_n_83));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b11___05F05d (.D(dbg_0_n_83),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[11]),.QN());
	NOR4_X1_LVT dbg_0i_37_2 (.A1(dbg_0_mem_cnt[8]),.A2(dbg_0_mem_cnt[9]),.A3(dbg_0_mem_cnt[10]),.A4(dbg_0_mem_cnt[11]),.ZN(dbg_0_n_37_2));
	OR2_X1_LVT dbg_0i_39_25 (.A1(dbg_0_mem_cnt[11]),.A2(dbg_0_n_39_12),.ZN(dbg_0_n_39_13));
	XNOR2_X1_LVT dbg_0i_39_26 (.A(dbg_0_mem_cnt[12]),.B(dbg_0_n_39_13),.ZN(dbg_0_n_68));
	AOI22_X1_LVT dbg_0i_40_25 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_68),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[12]),.ZN(dbg_0_n_40_13));
	INV_X1_LVT dbg_0i_40_26 (.A(dbg_0_n_40_13),.ZN(dbg_0_n_84));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b12___05F05d (.D(dbg_0_n_84),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[12]),.QN());
	OR2_X1_LVT dbg_0i_39_27 (.A1(dbg_0_mem_cnt[12]),.A2(dbg_0_n_39_13),.ZN(dbg_0_n_39_14));
	XNOR2_X1_LVT dbg_0i_39_28 (.A(dbg_0_mem_cnt[13]),.B(dbg_0_n_39_14),.ZN(dbg_0_n_69));
	AOI22_X1_LVT dbg_0i_40_27 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_69),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[13]),.ZN(dbg_0_n_40_14));
	INV_X1_LVT dbg_0i_40_28 (.A(dbg_0_n_40_14),.ZN(dbg_0_n_85));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b13___05F05d (.D(dbg_0_n_85),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[13]),.QN());
	OR2_X1_LVT dbg_0i_39_29 (.A1(dbg_0_mem_cnt[13]),.A2(dbg_0_n_39_14),.ZN(dbg_0_n_39_15));
	XNOR2_X1_LVT dbg_0i_39_30 (.A(dbg_0_mem_cnt[14]),.B(dbg_0_n_39_15),.ZN(dbg_0_n_70));
	AOI22_X1_LVT dbg_0i_40_29 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_70),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[14]),.ZN(dbg_0_n_40_15));
	INV_X1_LVT dbg_0i_40_30 (.A(dbg_0_n_40_15),.ZN(dbg_0_n_86));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b14___05F05d (.D(dbg_0_n_86),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[14]),.QN());
	OR2_X1_LVT dbg_0i_39_31 (.A1(dbg_0_mem_cnt[14]),.A2(dbg_0_n_39_15),.ZN(dbg_0_n_39_16));
	XNOR2_X1_LVT dbg_0i_39_32 (.A(dbg_0_mem_cnt[15]),.B(dbg_0_n_39_16),.ZN(dbg_0_n_71));
	AOI22_X1_LVT dbg_0i_40_31 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_71),.B1(dbg_0_n_102),.B2(dbg_0_dbg_din[15]),.ZN(dbg_0_n_40_16));
	INV_X1_LVT dbg_0i_40_32 (.A(dbg_0_n_40_16),.ZN(dbg_0_n_87));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b15___05F05d (.D(dbg_0_n_87),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[15]),.QN());
	NOR4_X1_LVT dbg_0i_37_3 (.A1(dbg_0_mem_cnt[12]),.A2(dbg_0_mem_cnt[13]),.A3(dbg_0_mem_cnt[14]),.A4(dbg_0_mem_cnt[15]),.ZN(dbg_0_n_37_3));
	NAND4_X1_LVT dbg_0i_37_4 (.A1(dbg_0_n_37_0),.A2(dbg_0_n_37_1),.A3(dbg_0_n_37_2),.A4(dbg_0_n_37_3),.ZN(dbg_0_n_37_4));
	CLKGATETST_X1_LVT dbg_0clk_gate_mem_ctl_reg (.CK(dbg_clk),.E(dbg_0_mem_ctl_wr),.SE(1'b0),.GCK(dbg_0_n_2));
	DFFR_X1_LVT dbg_0mem_ctl_reg___05F05b1___05F05d (.D(dbg_0_dbg_din[1]),.RN(dbg_0_n_104),.CK(dbg_0_n_2),.Q(dbg_0_mem_ctl[0]),.QN());
	OAI21_X1_LVT dbg_0i_6_0 (.A(dbg_0_mem_burst),.B1(dbg_0_dbg_wr),.B2(dbg_0_dbg_rd),.ZN(dbg_0_n_6_0));
	INV_X1_LVT dbg_0i_4_0 (.A(dbg_0_mem_ctl[0]),.ZN(dbg_0_n_3));
	AND2_X1_LVT dbg_0i_5_0 (.A1(dbg_0_n_3),.A2(dbg_0_mem_burst_start),.ZN(dbg_0_mem_burst_rd));
	INV_X1_LVT dbg_0i_6_1 (.A(dbg_0_mem_burst_rd),.ZN(dbg_0_n_6_1));
	NAND2_X1_LVT dbg_0i_6_2 (.A1(dbg_0_n_6_0),.A2(dbg_0_n_6_1),.ZN(dbg_0_n_4));
	DFFR_X1_LVT dbg_0mem_startb_reg (.D(dbg_0_n_4),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_startb),.QN());
	NOR4_X1_LVT dbg_0i_0_0 (.A1(dbg_0_mem_cnt[0]),.A2(dbg_0_mem_cnt[1]),.A3(dbg_0_mem_cnt[2]),.A4(dbg_0_mem_cnt[3]),.ZN(dbg_0_n_0_0));
	NOR4_X1_LVT dbg_0i_0_1 (.A1(dbg_0_mem_cnt[4]),.A2(dbg_0_mem_cnt[5]),.A3(dbg_0_mem_cnt[6]),.A4(dbg_0_mem_cnt[7]),.ZN(dbg_0_n_0_1));
	NOR4_X1_LVT dbg_0i_0_2 (.A1(dbg_0_mem_cnt[8]),.A2(dbg_0_mem_cnt[9]),.A3(dbg_0_mem_cnt[10]),.A4(dbg_0_mem_cnt[11]),.ZN(dbg_0_n_0_2));
	NOR4_X1_LVT dbg_0i_0_3 (.A1(dbg_0_mem_cnt[12]),.A2(dbg_0_mem_cnt[13]),.A3(dbg_0_mem_cnt[14]),.A4(dbg_0_mem_cnt[15]),.ZN(dbg_0_n_0_3));
	AND4_X1_LVT dbg_0i_0_4 (.A1(dbg_0_n_0_0),.A2(dbg_0_n_0_1),.A3(dbg_0_n_0_2),.A4(dbg_0_n_0_3),.ZN(dbg_0_n_0));
	AOI21_X1_LVT dbg_0i_8_0 (.A(dbg_0_mem_startb),.B1(dbg_0_n_0),.B2(dbg_0_mem_start),.ZN(dbg_0_n_8_0));
	INV_X1_LVT dbg_0i_8_1 (.A(dbg_0_n_8_0),.ZN(dbg_0_n_5));
	NAND2_X1_LVT dbg_0i_9_0 (.A1(cpu_halt_st),.A2(dbg_0_n_5),.ZN(dbg_0_n_9_0));
	INV_X1_LVT dbg_0i_9_1 (.A(dbg_0_n_9_0),.ZN(dbg_0_n_9_1));
	INV_X1_LVT dbg_0i_9_7 (.A(cpu_halt_st),.ZN(dbg_0_n_9_6));
	AOI21_X1_LVT dbg_0i_9_2 (.A(dbg_0_n_9_1),.B1(dbg_0_n_9_6),.B2(dbg_0_n_5),.ZN(dbg_0_n_9_2));
	INV_X1_LVT dbg_0i_9_4 (.A(dbg_0_mem_state[1]),.ZN(dbg_0_n_9_4));
	NAND2_X1_LVT dbg_0i_9_5 (.A1(dbg_0_n_9_4),.A2(dbg_0_mem_state[0]),.ZN(dbg_0_n_9_5));
	OAI22_X1_LVT dbg_0i_9_8 (.A1(dbg_0_n_9_3),.A2(dbg_0_n_9_0),.B1(dbg_0_n_9_5),.B2(dbg_0_n_9_6),.ZN(dbg_0_mem_state_nxt_reg[1]));
	DFFR_X1_LVT dbg_0mem_state_reg___05F05b1___05F05d (.D(dbg_0_mem_state_nxt_reg[1]),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_state[1]),.QN());
	OR2_X1_LVT dbg_0i_9_3 (.A1(dbg_0_mem_state[0]),.A2(dbg_0_mem_state[1]),.ZN(dbg_0_n_9_3));
	OAI22_X1_LVT dbg_0i_9_6 (.A1(dbg_0_n_9_2),.A2(dbg_0_n_9_3),.B1(dbg_0_n_9_5),.B2(cpu_halt_st),.ZN(dbg_0_mem_state_nxt_reg[0]));
	DFFR_X1_LVT dbg_0mem_state_reg___05F05b0___05F05d (.D(dbg_0_mem_state_nxt_reg[0]),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_state[0]),.QN());
	AND2_X1_LVT dbg_0i_12_0 (.A1(dbg_0_mem_state[0]),.A2(dbg_0_mem_state[1]),.ZN(dbg_0_n_6));
	INV_X1_LVT dbg_0i_12_1 (.A(dbg_0_mem_state[1]),.ZN(dbg_0_n_12_0));
	NOR2_X1_LVT dbg_0i_12_2 (.A1(dbg_0_n_12_0),.A2(dbg_0_mem_state[0]),.ZN(dbg_0_n_7));
	OR2_X1_LVT dbg_0i_13_0 (.A1(dbg_0_n_6),.A2(dbg_0_n_7),.ZN(dbg_0_mem_access));
	DFFR_X1_LVT dbg_0mem_ctl_reg___05F05b2___05F05d (.D(dbg_0_dbg_din[2]),.RN(dbg_0_n_104),.CK(dbg_0_n_2),.Q(dbg_0_mem_ctl[1]),.QN());
	INV_X1_LVT dbg_0i_23_0 (.A(dbg_0_mem_ctl[1]),.ZN(dbg_0_n_47));
	AND2_X1_LVT dbg_0i_24_0 (.A1(dbg_0_mem_access),.A2(dbg_0_n_47),.ZN(dbg_mem_en));
	AND2_X1_LVT dbg_0i_25_0 (.A1(dbg_0_mem_ctl[0]),.A2(dbg_mem_en),.ZN(dbg_0_n_48));
	NOR2_X1_LVT dbg_0i_49_3 (.A1(dbg_0_n_49_0),.A2(dbg_0_dbg_addr_in[1]),.ZN(dbg_0_n_49_3));
	NAND2_X1_LVT dbg_0i_49_12 (.A1(dbg_0_n_49_3),.A2(dbg_0_dbg_addr_in[2]),.ZN(dbg_0_n_49_12));
	NOR2_X1_LVT dbg_0i_49_27 (.A1(dbg_0_n_49_12),.A2(dbg_0_n_49_20),.ZN(dbg_0_n_96));
	AND2_X1_LVT dbg_0i_50_3 (.A1(dbg_0_dbg_wr),.A2(dbg_0_n_96),.ZN(dbg_0_n_101));
	INV_X1_LVT dbg_0i_20_0 (.A(dbg_0_n_101),.ZN(dbg_0_n_20_0));
	NOR4_X1_LVT dbg_0i_17_0 (.A1(dbg_0_mem_cnt[0]),.A2(dbg_0_mem_cnt[1]),.A3(dbg_0_mem_cnt[2]),.A4(dbg_0_mem_cnt[3]),.ZN(dbg_0_n_17_0));
	NOR4_X1_LVT dbg_0i_17_1 (.A1(dbg_0_mem_cnt[4]),.A2(dbg_0_mem_cnt[5]),.A3(dbg_0_mem_cnt[6]),.A4(dbg_0_mem_cnt[7]),.ZN(dbg_0_n_17_1));
	NOR4_X1_LVT dbg_0i_17_2 (.A1(dbg_0_mem_cnt[8]),.A2(dbg_0_mem_cnt[9]),.A3(dbg_0_mem_cnt[10]),.A4(dbg_0_mem_cnt[11]),.ZN(dbg_0_n_17_2));
	NOR4_X1_LVT dbg_0i_17_3 (.A1(dbg_0_mem_cnt[12]),.A2(dbg_0_mem_cnt[13]),.A3(dbg_0_mem_cnt[14]),.A4(dbg_0_mem_cnt[15]),.ZN(dbg_0_n_17_3));
	NAND4_X1_LVT dbg_0i_17_4 (.A1(dbg_0_n_17_0),.A2(dbg_0_n_17_1),.A3(dbg_0_n_17_2),.A4(dbg_0_n_17_3),.ZN(dbg_0_n_17_4));
	INV_X1_LVT dbg_0i_16_0 (.A(dbg_0_dbg_mem_acc),.ZN(dbg_0_n_16_0));
	DFFR_X1_LVT dbg_0mem_ctl_reg___05F05b3___05F05d (.D(dbg_0_dbg_din[3]),.RN(dbg_0_n_104),.CK(dbg_0_n_2),.Q(dbg_0_mem_ctl[2]),.QN());
	NOR2_X1_LVT dbg_0i_16_1 (.A1(dbg_0_n_16_0),.A2(dbg_0_mem_ctl[2]),.ZN(dbg_0_n_10));
	NAND2_X1_LVT dbg_0i_17_5 (.A1(dbg_0_n_10),.A2(dbg_0_mem_burst),.ZN(dbg_0_n_17_5));
	AND4_X1_LVT dbg_0i_17_6 (.A1(dbg_0_n_17_4),.A2(dbg_0_n_17_5),.A3(dbg_0_mem_burst),.A4(dbg_0_n_53),.ZN(dbg_0_n_11));
	HA_X1_LVT dbg_0i_19_0 (.A(dbg_0_n_11),.B(dbg_mem_addr[0]),.CO(dbg_0_n_19_0),.S(dbg_0_n_13));
	AOI22_X1_LVT dbg_0i_20_1 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_13),.B1(dbg_0_dbg_din[0]),.B2(dbg_0_n_101),.ZN(dbg_0_n_20_1));
	INV_X1_LVT dbg_0i_20_2 (.A(dbg_0_n_20_1),.ZN(dbg_0_n_29));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b0___05F05d (.D(dbg_0_n_29),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[0]),.QN());
	NAND2_X1_LVT dbg_0i_22_2 (.A1(dbg_mem_addr[0]),.A2(dbg_0_mem_ctl[2]),.ZN(dbg_0_n_46));
	AND2_X1_LVT dbg_0i_26_0 (.A1(dbg_0_n_48),.A2(dbg_0_n_46),.ZN(dbg_mem_wr[0]));
	INV_X1_LVT dbg_0i_22_0 (.A(dbg_mem_addr[0]),.ZN(dbg_0_n_22_0));
	NAND2_X1_LVT dbg_0i_22_1 (.A1(dbg_0_n_22_0),.A2(dbg_0_mem_ctl[2]),.ZN(dbg_0_n_45));
	AND2_X1_LVT dbg_0i_26_1 (.A1(dbg_0_n_48),.A2(dbg_0_n_45),.ZN(dbg_mem_wr[1]));
	OR2_X1_LVT dbg_0i_27_0 (.A1(dbg_mem_wr[0]),.A2(dbg_mem_wr[1]),.ZN(dbg_0_n_49));
	OR2_X1_LVT dbg_0i_31_0 (.A1(dbg_0_mem_burst),.A2(dbg_0_mem_burst_rd),.ZN(dbg_0_n_51));
	INV_X1_LVT dbg_0i_32_0 (.A(dbg_0_n_51),.ZN(dbg_0_n_32_0));
	AND2_X1_LVT dbg_0i_14_0 (.A1(dbg_0_mem_ctl[1]),.A2(dbg_0_mem_access),.ZN(dbg_0_n_9));
	AND2_X1_LVT dbg_0i_28_0 (.A1(dbg_0_n_3),.A2(dbg_0_n_9),.ZN(dbg_0_dbg_reg_rd));
	AND2_X1_LVT dbg_0i_29_0 (.A1(dbg_0_n_3),.A2(dbg_mem_en),.ZN(dbg_0_dbg_mem_rd));
	DFFR_X1_LVT dbg_0dbg_mem_rd_dly_reg (.D(dbg_0_dbg_mem_rd),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_dbg_mem_rd_dly),.QN());
	OR2_X1_LVT dbg_0i_30_0 (.A1(dbg_0_dbg_reg_rd),.A2(dbg_0_dbg_mem_rd_dly),.ZN(dbg_0_n_50));
	AOI22_X1_LVT dbg_0i_32_1 (.A1(dbg_0_n_32_0),.A2(dbg_0_dbg_rd),.B1(dbg_0_n_50),.B2(dbg_0_n_51),.ZN(dbg_0_n_32_1));
	INV_X1_LVT dbg_0i_32_2 (.A(dbg_0_n_32_1),.ZN(dbg_0_n_52));
	DFFR_X1_LVT dbg_0dbg_rd_rdy_reg (.D(dbg_0_n_52),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_dbg_rd_rdy),.QN());
	AOI21_X1_LVT dbg_0i_34_0 (.A(dbg_0_n_49),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_n_47),.ZN(dbg_0_n_34_0));
	INV_X1_LVT dbg_0i_34_1 (.A(dbg_0_n_34_0),.ZN(dbg_0_dbg_mem_acc));
	AND2_X1_LVT dbg_0i_15_0 (.A1(dbg_0_mem_ctl[0]),.A2(dbg_0_n_9),.ZN(dbg_reg_wr));
	NOR2_X1_LVT dbg_0i_35_0 (.A1(dbg_0_dbg_mem_acc),.A2(dbg_reg_wr),.ZN(dbg_0_n_35_0));
	NAND2_X1_LVT dbg_0i_35_1 (.A1(dbg_0_mem_ctl[1]),.A2(dbg_0_dbg_rd_rdy),.ZN(dbg_0_n_35_1));
	NAND2_X1_LVT dbg_0i_35_2 (.A1(dbg_0_n_35_0),.A2(dbg_0_n_35_1),.ZN(dbg_0_n_53));
	AND2_X1_LVT dbg_0i_36_0 (.A1(dbg_0_n_53),.A2(dbg_0_mem_burst),.ZN(dbg_0_n_54));
	AND2_X1_LVT dbg_0i_37_5 (.A1(dbg_0_n_37_4),.A2(dbg_0_n_54),.ZN(dbg_0_n_55));
	XNOR2_X1_LVT dbg_0i_39_0 (.A(dbg_0_n_55),.B(dbg_0_mem_cnt[0]),.ZN(dbg_0_n_39_0));
	INV_X1_LVT dbg_0i_39_1 (.A(dbg_0_n_39_0),.ZN(dbg_0_n_56));
	AOI22_X1_LVT dbg_0i_40_1 (.A1(dbg_0_n_40_0),.A2(dbg_0_n_56),.B1(dbg_0_dbg_din[0]),.B2(dbg_0_n_102),.ZN(dbg_0_n_40_1));
	INV_X1_LVT dbg_0i_40_2 (.A(dbg_0_n_40_1),.ZN(dbg_0_n_72));
	DFFR_X1_LVT dbg_0mem_cnt_reg___05F05b0___05F05d (.D(dbg_0_n_72),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_mem_cnt[0]),.QN());
	NOR4_X1_LVT dbg_0i_42_0 (.A1(dbg_0_mem_cnt[0]),.A2(dbg_0_mem_cnt[1]),.A3(dbg_0_mem_cnt[2]),.A4(dbg_0_mem_cnt[3]),.ZN(dbg_0_n_42_0));
	NOR4_X1_LVT dbg_0i_42_1 (.A1(dbg_0_mem_cnt[4]),.A2(dbg_0_mem_cnt[5]),.A3(dbg_0_mem_cnt[6]),.A4(dbg_0_mem_cnt[7]),.ZN(dbg_0_n_42_1));
	NOR4_X1_LVT dbg_0i_42_2 (.A1(dbg_0_mem_cnt[8]),.A2(dbg_0_mem_cnt[9]),.A3(dbg_0_mem_cnt[10]),.A4(dbg_0_mem_cnt[11]),.ZN(dbg_0_n_42_2));
	NOR4_X1_LVT dbg_0i_42_3 (.A1(dbg_0_mem_cnt[12]),.A2(dbg_0_mem_cnt[13]),.A3(dbg_0_mem_cnt[14]),.A4(dbg_0_mem_cnt[15]),.ZN(dbg_0_n_42_3));
	NAND4_X1_LVT dbg_0i_42_4 (.A1(dbg_0_n_42_0),.A2(dbg_0_n_42_1),.A3(dbg_0_n_42_2),.A4(dbg_0_n_42_3),.ZN(dbg_0_n_88));
	AND2_X1_LVT dbg_0i_43_0 (.A1(dbg_0_mem_start),.A2(dbg_0_n_88),.ZN(dbg_0_mem_burst_start));
	OAI21_X1_LVT dbg_0i_44_0 (.A(dbg_0_n_0),.B1(dbg_0_dbg_wr),.B2(dbg_0_dbg_rd_rdy),.ZN(dbg_0_n_44_0));
	INV_X1_LVT dbg_0i_44_1 (.A(dbg_0_n_44_0),.ZN(dbg_0_mem_burst_end));
	INV_X1_LVT dbg_0i_46_1 (.A(dbg_0_mem_burst_end),.ZN(dbg_0_n_46_1));
	INV_X1_LVT dbg_0i_46_0 (.A(dbg_0_mem_burst_start),.ZN(dbg_0_n_46_0));
	NAND2_X1_LVT dbg_0i_46_2 (.A1(dbg_0_n_46_1),.A2(dbg_0_n_46_0),.ZN(dbg_0_n_90));
	CLKGATETST_X1_LVT dbg_0clk_gate_mem_burst_reg (.CK(dbg_clk),.E(dbg_0_n_90),.SE(1'b0),.GCK(dbg_0_n_89));
	DFFR_X1_LVT dbg_0mem_burst_reg (.D(dbg_0_mem_burst_start),.RN(dbg_0_n_104),.CK(dbg_0_n_89),.Q(dbg_0_mem_burst),.QN());
	INV_X1_LVT dbg_0i_48_0 (.A(dbg_0_mem_burst),.ZN(dbg_0_n_48_0));
	AND2_X1_LVT dbg_0i_48_1 (.A1(dbg_0_n_48_0),.A2(dbg_0_dbg_addr[0]),.ZN(dbg_0_dbg_addr_in[0]));
	INV_X1_LVT dbg_0i_49_0 (.A(dbg_0_dbg_addr_in[0]),.ZN(dbg_0_n_49_0));
	INV_X1_LVT dbg_0i_49_1 (.A(dbg_0_dbg_addr_in[1]),.ZN(dbg_0_n_49_1));
	NOR2_X1_LVT dbg_0i_49_5 (.A1(dbg_0_n_49_0),.A2(dbg_0_n_49_1),.ZN(dbg_0_n_49_5));
	NAND2_X1_LVT dbg_0i_49_14 (.A1(dbg_0_n_49_5),.A2(dbg_0_dbg_addr_in[2]),.ZN(dbg_0_n_49_14));
	NOR2_X1_LVT dbg_0i_49_29 (.A1(dbg_0_n_49_14),.A2(dbg_0_n_49_20),.ZN(dbg_0_n_98));
	NAND2_X1_LVT dbg_0i_78_125 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[15]),.ZN(dbg_0_n_78_110));
	AOI22_X1_LVT dbg_0i_20_29 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_27),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[14]),.ZN(dbg_0_n_20_15));
	INV_X1_LVT dbg_0i_20_30 (.A(dbg_0_n_20_15),.ZN(dbg_0_n_43));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b14___05F05d (.D(dbg_0_n_43),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[14]),.QN());
	AOI22_X1_LVT dbg_0i_20_27 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_26),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[13]),.ZN(dbg_0_n_20_14));
	INV_X1_LVT dbg_0i_20_28 (.A(dbg_0_n_20_14),.ZN(dbg_0_n_42));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b13___05F05d (.D(dbg_0_n_42),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[13]),.QN());
	AOI22_X1_LVT dbg_0i_20_25 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_25),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[12]),.ZN(dbg_0_n_20_13));
	INV_X1_LVT dbg_0i_20_26 (.A(dbg_0_n_20_13),.ZN(dbg_0_n_41));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b12___05F05d (.D(dbg_0_n_41),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[12]),.QN());
	AOI22_X1_LVT dbg_0i_20_23 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_24),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[11]),.ZN(dbg_0_n_20_12));
	INV_X1_LVT dbg_0i_20_24 (.A(dbg_0_n_20_12),.ZN(dbg_0_n_40));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b11___05F05d (.D(dbg_0_n_40),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[11]),.QN());
	AOI22_X1_LVT dbg_0i_20_21 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_23),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[10]),.ZN(dbg_0_n_20_11));
	INV_X1_LVT dbg_0i_20_22 (.A(dbg_0_n_20_11),.ZN(dbg_0_n_39));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b10___05F05d (.D(dbg_0_n_39),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[10]),.QN());
	AOI22_X1_LVT dbg_0i_20_19 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_22),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[9]),.ZN(dbg_0_n_20_10));
	INV_X1_LVT dbg_0i_20_20 (.A(dbg_0_n_20_10),.ZN(dbg_0_n_38));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b9___05F05d (.D(dbg_0_n_38),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[9]),.QN());
	AOI22_X1_LVT dbg_0i_20_17 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_21),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[8]),.ZN(dbg_0_n_20_9));
	INV_X1_LVT dbg_0i_20_18 (.A(dbg_0_n_20_9),.ZN(dbg_0_n_37));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b8___05F05d (.D(dbg_0_n_37),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[8]),.QN());
	AOI22_X1_LVT dbg_0i_20_15 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_20),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[7]),.ZN(dbg_0_n_20_8));
	INV_X1_LVT dbg_0i_20_16 (.A(dbg_0_n_20_8),.ZN(dbg_0_n_36));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b7___05F05d (.D(dbg_0_n_36),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[7]),.QN());
	AOI22_X1_LVT dbg_0i_20_13 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_19),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[6]),.ZN(dbg_0_n_20_7));
	INV_X1_LVT dbg_0i_20_14 (.A(dbg_0_n_20_7),.ZN(dbg_0_n_35));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b6___05F05d (.D(dbg_0_n_35),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[6]),.QN());
	AOI22_X1_LVT dbg_0i_20_11 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_18),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[5]),.ZN(dbg_0_n_20_6));
	INV_X1_LVT dbg_0i_20_12 (.A(dbg_0_n_20_6),.ZN(dbg_0_n_34));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b5___05F05d (.D(dbg_0_n_34),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[5]),.QN());
	AOI22_X1_LVT dbg_0i_20_9 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_17),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[4]),.ZN(dbg_0_n_20_5));
	INV_X1_LVT dbg_0i_20_10 (.A(dbg_0_n_20_5),.ZN(dbg_0_n_33));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b4___05F05d (.D(dbg_0_n_33),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[4]),.QN());
	AOI22_X1_LVT dbg_0i_20_7 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_16),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[3]),.ZN(dbg_0_n_20_4));
	INV_X1_LVT dbg_0i_20_8 (.A(dbg_0_n_20_4),.ZN(dbg_0_n_32));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b3___05F05d (.D(dbg_0_n_32),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[3]),.QN());
	AOI22_X1_LVT dbg_0i_20_5 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_15),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[2]),.ZN(dbg_0_n_20_3));
	INV_X1_LVT dbg_0i_20_6 (.A(dbg_0_n_20_3),.ZN(dbg_0_n_31));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b2___05F05d (.D(dbg_0_n_31),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[2]),.QN());
	INV_X1_LVT dbg_0i_17_7 (.A(dbg_0_n_17_4),.ZN(dbg_0_n_17_6));
	NOR2_X1_LVT dbg_0i_17_8 (.A1(dbg_0_n_17_6),.A2(dbg_0_n_17_5),.ZN(dbg_0_n_12));
	AOI22_X1_LVT dbg_0i_20_3 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_14),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[1]),.ZN(dbg_0_n_20_2));
	INV_X1_LVT dbg_0i_20_4 (.A(dbg_0_n_20_2),.ZN(dbg_0_n_30));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b1___05F05d (.D(dbg_0_n_30),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[1]),.QN());
	FA_X1_LVT dbg_0i_19_1 (.A(dbg_0_n_12),.B(dbg_mem_addr[1]),.CI(dbg_0_n_19_0),.CO(dbg_0_n_19_1),.S(dbg_0_n_14));
	HA_X1_LVT dbg_0i_19_2 (.A(dbg_mem_addr[2]),.B(dbg_0_n_19_1),.CO(dbg_0_n_19_2),.S(dbg_0_n_15));
	HA_X1_LVT dbg_0i_19_3 (.A(dbg_mem_addr[3]),.B(dbg_0_n_19_2),.CO(dbg_0_n_19_3),.S(dbg_0_n_16));
	HA_X1_LVT dbg_0i_19_4 (.A(dbg_mem_addr[4]),.B(dbg_0_n_19_3),.CO(dbg_0_n_19_4),.S(dbg_0_n_17));
	HA_X1_LVT dbg_0i_19_5 (.A(dbg_mem_addr[5]),.B(dbg_0_n_19_4),.CO(dbg_0_n_19_5),.S(dbg_0_n_18));
	HA_X1_LVT dbg_0i_19_6 (.A(dbg_mem_addr[6]),.B(dbg_0_n_19_5),.CO(dbg_0_n_19_6),.S(dbg_0_n_19));
	HA_X1_LVT dbg_0i_19_7 (.A(dbg_mem_addr[7]),.B(dbg_0_n_19_6),.CO(dbg_0_n_19_7),.S(dbg_0_n_20));
	HA_X1_LVT dbg_0i_19_8 (.A(dbg_mem_addr[8]),.B(dbg_0_n_19_7),.CO(dbg_0_n_19_8),.S(dbg_0_n_21));
	HA_X1_LVT dbg_0i_19_9 (.A(dbg_mem_addr[9]),.B(dbg_0_n_19_8),.CO(dbg_0_n_19_9),.S(dbg_0_n_22));
	HA_X1_LVT dbg_0i_19_10 (.A(dbg_mem_addr[10]),.B(dbg_0_n_19_9),.CO(dbg_0_n_19_10),.S(dbg_0_n_23));
	HA_X1_LVT dbg_0i_19_11 (.A(dbg_mem_addr[11]),.B(dbg_0_n_19_10),.CO(dbg_0_n_19_11),.S(dbg_0_n_24));
	HA_X1_LVT dbg_0i_19_12 (.A(dbg_mem_addr[12]),.B(dbg_0_n_19_11),.CO(dbg_0_n_19_12),.S(dbg_0_n_25));
	HA_X1_LVT dbg_0i_19_13 (.A(dbg_mem_addr[13]),.B(dbg_0_n_19_12),.CO(dbg_0_n_19_13),.S(dbg_0_n_26));
	HA_X1_LVT dbg_0i_19_14 (.A(dbg_mem_addr[14]),.B(dbg_0_n_19_13),.CO(dbg_0_n_19_14),.S(dbg_0_n_27));
	XNOR2_X1_LVT dbg_0i_19_15 (.A(dbg_mem_addr[15]),.B(dbg_0_n_19_14),.ZN(dbg_0_n_19_15));
	INV_X1_LVT dbg_0i_19_16 (.A(dbg_0_n_19_15),.ZN(dbg_0_n_28));
	AOI22_X1_LVT dbg_0i_20_31 (.A1(dbg_0_n_20_0),.A2(dbg_0_n_28),.B1(dbg_0_n_101),.B2(dbg_0_dbg_din[15]),.ZN(dbg_0_n_20_16));
	INV_X1_LVT dbg_0i_20_32 (.A(dbg_0_n_20_16),.ZN(dbg_0_n_44));
	DFFR_X1_LVT dbg_0mem_addr_reg___05F05b15___05F05d (.D(dbg_0_n_44),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_mem_addr[15]),.QN());
	NAND2_X1_LVT dbg_0i_78_126 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[15]),.ZN(dbg_0_n_78_111));
	NOR2_X1_LVT dbg_0i_49_4 (.A1(dbg_0_dbg_addr_in[0]),.A2(dbg_0_n_49_1),.ZN(dbg_0_n_49_4));
	NAND2_X1_LVT dbg_0i_49_13 (.A1(dbg_0_n_49_4),.A2(dbg_0_dbg_addr_in[2]),.ZN(dbg_0_n_49_13));
	NOR2_X1_LVT dbg_0i_49_28 (.A1(dbg_0_n_49_13),.A2(dbg_0_n_49_20),.ZN(dbg_0_n_97));
	AND2_X1_LVT dbg_0i_50_4 (.A1(dbg_0_dbg_wr),.A2(dbg_0_n_97),.ZN(dbg_0_mem_data_wr));
	INV_X1_LVT dbg_0i_70_1 (.A(dbg_0_dbg_reg_rd),.ZN(dbg_0_n_70_0));
	NOR2_X1_LVT dbg_0i_70_2 (.A1(dbg_0_n_70_0),.A2(dbg_0_mem_data_wr),.ZN(dbg_0_n_136));
	NOR2_X1_LVT dbg_0i_70_0 (.A1(dbg_0_dbg_reg_rd),.A2(dbg_0_mem_data_wr),.ZN(dbg_0_n_135));
	INV_X1_LVT dbg_0i_67_0 (.A(dbg_0_mem_ctl[2]),.ZN(dbg_0_n_115));
	AND2_X1_LVT dbg_0i_68_24 (.A1(dbg_0_n_115),.A2(dbg_mem_din[15]),.ZN(dbg_0_n_133));
	AOI222_X1_LVT dbg_0i_71_30 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[15]),.B1(dbg_0_n_136),.B2(dbg_reg_din[15]),.C1(dbg_0_n_135),.C2(dbg_0_n_133),.ZN(dbg_0_n_71_15));
	INV_X1_LVT dbg_0i_71_31 (.A(dbg_0_n_71_15),.ZN(dbg_0_n_152));
	INV_X1_LVT dbg_0i_72_0 (.A(dbg_0_dbg_reg_rd),.ZN(dbg_0_n_72_0));
	INV_X1_LVT dbg_0i_72_1 (.A(dbg_0_mem_data_wr),.ZN(dbg_0_n_72_1));
	NAND3_X1_LVT dbg_0i_72_2 (.A1(dbg_0_n_72_0),.A2(dbg_0_n_72_1),.A3(dbg_0_dbg_mem_rd_dly),.ZN(dbg_0_n_72_2));
	NAND3_X1_LVT dbg_0i_72_3 (.A1(dbg_0_n_72_2),.A2(dbg_0_n_72_0),.A3(dbg_0_n_72_1),.ZN(dbg_0_n_153));
	CLKGATETST_X1_LVT dbg_0clk_gate_mem_data_reg (.CK(dbg_clk),.E(dbg_0_n_153),.SE(1'b0),.GCK(dbg_0_n_134));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b15___05F05d (.D(dbg_0_n_152),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[15]),.QN());
	NAND2_X1_LVT dbg_0i_78_127 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[15]),.ZN(dbg_0_n_78_112));
	INV_X1_LVT dbg_0i_49_6 (.A(dbg_0_dbg_addr_in[2]),.ZN(dbg_0_n_49_6));
	NAND2_X1_LVT dbg_0i_49_8 (.A1(dbg_0_n_49_3),.A2(dbg_0_n_49_6),.ZN(dbg_0_n_49_8));
	NOR2_X1_LVT dbg_0i_49_23 (.A1(dbg_0_n_49_8),.A2(dbg_0_n_49_20),.ZN(dbg_0_n_92));
	NAND2_X1_LVT dbg_0i_78_128 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_113));
	NAND4_X1_LVT dbg_0i_78_129 (.A1(dbg_0_n_78_110),.A2(dbg_0_n_78_111),.A3(dbg_0_n_78_112),.A4(dbg_0_n_78_113),.ZN(dbg_0_n_78_114));
	NAND2_X1_LVT dbg_0i_49_7 (.A1(dbg_0_n_49_2),.A2(dbg_0_n_49_6),.ZN(dbg_0_n_49_7));
	NOR2_X1_LVT dbg_0i_49_22 (.A1(dbg_0_n_49_7),.A2(dbg_0_n_49_20),.ZN(dbg_0_n_91));
	INV_X1_LVT dbg_0i_49_18 (.A(dbg_0_dbg_addr_in[5]),.ZN(dbg_0_n_49_18));
	NAND2_X1_LVT dbg_0i_49_17 (.A1(dbg_0_dbg_addr_in[4]),.A2(dbg_0_n_49_18),.ZN(dbg_0_n_49_17));
	INV_X1_LVT dbg_0i_49_19 (.A(dbg_0_n_49_17),.ZN(dbg_0_n_49_19));
	NAND2_X1_LVT dbg_0i_49_21 (.A1(dbg_0_dbg_addr_in[3]),.A2(dbg_0_n_49_19),.ZN(dbg_0_n_49_21));
	NOR2_X1_LVT dbg_0i_49_30 (.A1(dbg_0_n_49_7),.A2(dbg_0_n_49_21),.ZN(dbg_0_n_99));
	AOI221_X1_LVT dbg_0i_78_130 (.A(dbg_0_n_78_114),.B1(dbg_0_n_91),.B2(cpu_id[15]),.C1(dbg_0_n_99),.C2(1'b0),.ZN(dbg_0_n_78_115));
	INV_X1_LVT dbg_0i_78_131 (.A(dbg_0_n_78_115),.ZN(dbg_0_dbg_dout[15]));
	NAND2_X1_LVT dbg_0i_78_118 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[14]),.ZN(dbg_0_n_78_104));
	NAND2_X1_LVT dbg_0i_78_119 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[14]),.ZN(dbg_0_n_78_105));
	AND2_X1_LVT dbg_0i_68_23 (.A1(dbg_0_n_115),.A2(dbg_mem_din[14]),.ZN(dbg_0_n_132));
	AOI222_X1_LVT dbg_0i_71_28 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[14]),.B1(dbg_0_n_136),.B2(dbg_reg_din[14]),.C1(dbg_0_n_135),.C2(dbg_0_n_132),.ZN(dbg_0_n_71_14));
	INV_X1_LVT dbg_0i_71_29 (.A(dbg_0_n_71_14),.ZN(dbg_0_n_151));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b14___05F05d (.D(dbg_0_n_151),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[14]),.QN());
	NAND2_X1_LVT dbg_0i_78_120 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[14]),.ZN(dbg_0_n_78_106));
	NAND2_X1_LVT dbg_0i_78_121 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_107));
	NAND4_X1_LVT dbg_0i_78_122 (.A1(dbg_0_n_78_104),.A2(dbg_0_n_78_105),.A3(dbg_0_n_78_106),.A4(dbg_0_n_78_107),.ZN(dbg_0_n_78_108));
	AOI221_X1_LVT dbg_0i_78_123 (.A(dbg_0_n_78_108),.B1(dbg_0_n_91),.B2(cpu_id[14]),.C1(dbg_0_n_99),.C2(1'b0),.ZN(dbg_0_n_78_109));
	INV_X1_LVT dbg_0i_78_124 (.A(dbg_0_n_78_109),.ZN(dbg_0_dbg_dout[14]));
	NAND2_X1_LVT dbg_0i_78_111 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[13]),.ZN(dbg_0_n_78_98));
	NAND2_X1_LVT dbg_0i_78_112 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[13]),.ZN(dbg_0_n_78_99));
	AND2_X1_LVT dbg_0i_68_22 (.A1(dbg_0_n_115),.A2(dbg_mem_din[13]),.ZN(dbg_0_n_131));
	AOI222_X1_LVT dbg_0i_71_26 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[13]),.B1(dbg_0_n_136),.B2(dbg_reg_din[13]),.C1(dbg_0_n_135),.C2(dbg_0_n_131),.ZN(dbg_0_n_71_13));
	INV_X1_LVT dbg_0i_71_27 (.A(dbg_0_n_71_13),.ZN(dbg_0_n_150));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b13___05F05d (.D(dbg_0_n_150),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[13]),.QN());
	NAND2_X1_LVT dbg_0i_78_113 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[13]),.ZN(dbg_0_n_78_100));
	NAND2_X1_LVT dbg_0i_78_114 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_101));
	NAND4_X1_LVT dbg_0i_78_115 (.A1(dbg_0_n_78_98),.A2(dbg_0_n_78_99),.A3(dbg_0_n_78_100),.A4(dbg_0_n_78_101),.ZN(dbg_0_n_78_102));
	AOI221_X1_LVT dbg_0i_78_116 (.A(dbg_0_n_78_102),.B1(dbg_0_n_91),.B2(cpu_id[13]),.C1(dbg_0_n_99),.C2(1'b0),.ZN(dbg_0_n_78_103));
	INV_X1_LVT dbg_0i_78_117 (.A(dbg_0_n_78_103),.ZN(dbg_0_dbg_dout[13]));
	NAND2_X1_LVT dbg_0i_78_104 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[12]),.ZN(dbg_0_n_78_92));
	NAND2_X1_LVT dbg_0i_78_105 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[12]),.ZN(dbg_0_n_78_93));
	AND2_X1_LVT dbg_0i_68_21 (.A1(dbg_0_n_115),.A2(dbg_mem_din[12]),.ZN(dbg_0_n_130));
	AOI222_X1_LVT dbg_0i_71_24 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[12]),.B1(dbg_0_n_136),.B2(dbg_reg_din[12]),.C1(dbg_0_n_135),.C2(dbg_0_n_130),.ZN(dbg_0_n_71_12));
	INV_X1_LVT dbg_0i_71_25 (.A(dbg_0_n_71_12),.ZN(dbg_0_n_149));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b12___05F05d (.D(dbg_0_n_149),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[12]),.QN());
	NAND2_X1_LVT dbg_0i_78_106 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[12]),.ZN(dbg_0_n_78_94));
	NAND2_X1_LVT dbg_0i_78_107 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_95));
	NAND4_X1_LVT dbg_0i_78_108 (.A1(dbg_0_n_78_92),.A2(dbg_0_n_78_93),.A3(dbg_0_n_78_94),.A4(dbg_0_n_78_95),.ZN(dbg_0_n_78_96));
	AOI221_X1_LVT dbg_0i_78_109 (.A(dbg_0_n_78_96),.B1(dbg_0_n_91),.B2(cpu_id[12]),.C1(dbg_0_n_99),.C2(1'b0),.ZN(dbg_0_n_78_97));
	INV_X1_LVT dbg_0i_78_110 (.A(dbg_0_n_78_97),.ZN(dbg_0_dbg_dout[12]));
	NAND2_X1_LVT dbg_0i_78_97 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[11]),.ZN(dbg_0_n_78_86));
	NAND2_X1_LVT dbg_0i_78_98 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[11]),.ZN(dbg_0_n_78_87));
	AND2_X1_LVT dbg_0i_68_20 (.A1(dbg_0_n_115),.A2(dbg_mem_din[11]),.ZN(dbg_0_n_129));
	AOI222_X1_LVT dbg_0i_71_22 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[11]),.B1(dbg_0_n_136),.B2(dbg_reg_din[11]),.C1(dbg_0_n_135),.C2(dbg_0_n_129),.ZN(dbg_0_n_71_11));
	INV_X1_LVT dbg_0i_71_23 (.A(dbg_0_n_71_11),.ZN(dbg_0_n_148));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b11___05F05d (.D(dbg_0_n_148),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[11]),.QN());
	NAND2_X1_LVT dbg_0i_78_99 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[11]),.ZN(dbg_0_n_78_88));
	NAND2_X1_LVT dbg_0i_78_100 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_89));
	NAND4_X1_LVT dbg_0i_78_101 (.A1(dbg_0_n_78_86),.A2(dbg_0_n_78_87),.A3(dbg_0_n_78_88),.A4(dbg_0_n_78_89),.ZN(dbg_0_n_78_90));
	AOI221_X1_LVT dbg_0i_78_102 (.A(dbg_0_n_78_90),.B1(dbg_0_n_91),.B2(cpu_id[11]),.C1(dbg_0_n_99),.C2(1'b0),.ZN(dbg_0_n_78_91));
	INV_X1_LVT dbg_0i_78_103 (.A(dbg_0_n_78_91),.ZN(dbg_0_dbg_dout[11]));
	NAND2_X1_LVT dbg_0i_78_90 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[10]),.ZN(dbg_0_n_78_80));
	NAND2_X1_LVT dbg_0i_78_91 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[10]),.ZN(dbg_0_n_78_81));
	AND2_X1_LVT dbg_0i_68_19 (.A1(dbg_0_n_115),.A2(dbg_mem_din[10]),.ZN(dbg_0_n_128));
	AOI222_X1_LVT dbg_0i_71_20 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[10]),.B1(dbg_0_n_136),.B2(dbg_reg_din[10]),.C1(dbg_0_n_135),.C2(dbg_0_n_128),.ZN(dbg_0_n_71_10));
	INV_X1_LVT dbg_0i_71_21 (.A(dbg_0_n_71_10),.ZN(dbg_0_n_147));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b10___05F05d (.D(dbg_0_n_147),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[10]),.QN());
	NAND2_X1_LVT dbg_0i_78_92 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[10]),.ZN(dbg_0_n_78_82));
	NAND2_X1_LVT dbg_0i_78_93 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_83));
	NAND4_X1_LVT dbg_0i_78_94 (.A1(dbg_0_n_78_80),.A2(dbg_0_n_78_81),.A3(dbg_0_n_78_82),.A4(dbg_0_n_78_83),.ZN(dbg_0_n_78_84));
	AOI221_X1_LVT dbg_0i_78_95 (.A(dbg_0_n_78_84),.B1(dbg_0_n_91),.B2(cpu_id[10]),.C1(dbg_0_n_99),.C2(1'b0),.ZN(dbg_0_n_78_85));
	INV_X1_LVT dbg_0i_78_96 (.A(dbg_0_n_78_85),.ZN(dbg_0_dbg_dout[10]));
	NAND2_X1_LVT dbg_0i_78_83 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[9]),.ZN(dbg_0_n_78_74));
	NAND2_X1_LVT dbg_0i_78_84 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[9]),.ZN(dbg_0_n_78_75));
	AND2_X1_LVT dbg_0i_68_18 (.A1(dbg_0_n_115),.A2(dbg_mem_din[9]),.ZN(dbg_0_n_127));
	AOI222_X1_LVT dbg_0i_71_18 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[9]),.B1(dbg_0_n_136),.B2(dbg_reg_din[9]),.C1(dbg_0_n_135),.C2(dbg_0_n_127),.ZN(dbg_0_n_71_9));
	INV_X1_LVT dbg_0i_71_19 (.A(dbg_0_n_71_9),.ZN(dbg_0_n_146));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b9___05F05d (.D(dbg_0_n_146),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[9]),.QN());
	NAND2_X1_LVT dbg_0i_78_85 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[9]),.ZN(dbg_0_n_78_76));
	NAND2_X1_LVT dbg_0i_78_86 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_77));
	NAND4_X1_LVT dbg_0i_78_87 (.A1(dbg_0_n_78_74),.A2(dbg_0_n_78_75),.A3(dbg_0_n_78_76),.A4(dbg_0_n_78_77),.ZN(dbg_0_n_78_78));
	AOI221_X1_LVT dbg_0i_78_88 (.A(dbg_0_n_78_78),.B1(dbg_0_n_91),.B2(cpu_id[9]),.C1(dbg_0_n_99),.C2(1'b0),.ZN(dbg_0_n_78_79));
	INV_X1_LVT dbg_0i_78_89 (.A(dbg_0_n_78_79),.ZN(dbg_0_dbg_dout[9]));
	NAND2_X1_LVT dbg_0i_78_76 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[8]),.ZN(dbg_0_n_78_68));
	NAND2_X1_LVT dbg_0i_78_77 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[8]),.ZN(dbg_0_n_78_69));
	AND2_X1_LVT dbg_0i_68_17 (.A1(dbg_mem_din[8]),.A2(dbg_0_n_115),.ZN(dbg_0_n_126));
	AOI222_X1_LVT dbg_0i_71_16 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[8]),.B1(dbg_0_n_136),.B2(dbg_reg_din[8]),.C1(dbg_0_n_135),.C2(dbg_0_n_126),.ZN(dbg_0_n_71_8));
	INV_X1_LVT dbg_0i_71_17 (.A(dbg_0_n_71_8),.ZN(dbg_0_n_145));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b8___05F05d (.D(dbg_0_n_145),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[8]),.QN());
	NAND2_X1_LVT dbg_0i_78_78 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[8]),.ZN(dbg_0_n_78_70));
	NAND2_X1_LVT dbg_0i_78_79 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_71));
	NAND4_X1_LVT dbg_0i_78_80 (.A1(dbg_0_n_78_68),.A2(dbg_0_n_78_69),.A3(dbg_0_n_78_70),.A4(dbg_0_n_78_71),.ZN(dbg_0_n_78_72));
	AOI221_X1_LVT dbg_0i_78_81 (.A(dbg_0_n_78_72),.B1(dbg_0_n_91),.B2(cpu_id[8]),.C1(dbg_0_n_99),.C2(1'b0),.ZN(dbg_0_n_78_73));
	INV_X1_LVT dbg_0i_78_82 (.A(dbg_0_n_78_73),.ZN(dbg_0_dbg_dout[8]));
	NAND2_X1_LVT dbg_0i_78_69 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[7]),.ZN(dbg_0_n_78_62));
	NAND2_X1_LVT dbg_0i_78_70 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[7]),.ZN(dbg_0_n_78_63));
	NOR2_X1_LVT dbg_0i_67_1 (.A1(dbg_0_n_115),.A2(dbg_mem_addr[0]),.ZN(dbg_0_n_116));
	OR2_X1_LVT dbg_0i_68_0 (.A1(dbg_0_n_115),.A2(dbg_0_n_116),.ZN(dbg_0_n_68_0));
	AND2_X1_LVT dbg_0i_67_2 (.A1(dbg_mem_addr[0]),.A2(dbg_0_mem_ctl[2]),.ZN(dbg_0_n_117));
	AOI22_X1_LVT dbg_0i_68_15 (.A1(dbg_0_n_68_0),.A2(dbg_mem_din[7]),.B1(dbg_0_n_117),.B2(dbg_mem_din[15]),.ZN(dbg_0_n_68_8));
	INV_X1_LVT dbg_0i_68_16 (.A(dbg_0_n_68_8),.ZN(dbg_0_n_125));
	AOI222_X1_LVT dbg_0i_71_14 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[7]),.B1(dbg_0_n_136),.B2(dbg_reg_din[7]),.C1(dbg_0_n_135),.C2(dbg_0_n_125),.ZN(dbg_0_n_71_7));
	INV_X1_LVT dbg_0i_71_15 (.A(dbg_0_n_71_7),.ZN(dbg_0_n_144));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b7___05F05d (.D(dbg_0_n_144),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[7]),.QN());
	NAND2_X1_LVT dbg_0i_78_71 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[7]),.ZN(dbg_0_n_78_64));
	NAND2_X1_LVT dbg_0i_78_72 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_65));
	NAND4_X1_LVT dbg_0i_78_73 (.A1(dbg_0_n_78_62),.A2(dbg_0_n_78_63),.A3(dbg_0_n_78_64),.A4(dbg_0_n_78_65),.ZN(dbg_0_n_78_66));
	AOI221_X1_LVT dbg_0i_78_74 (.A(dbg_0_n_78_66),.B1(dbg_0_n_91),.B2(cpu_id[7]),.C1(dbg_0_n_99),.C2(1'b0),.ZN(dbg_0_n_78_67));
	INV_X1_LVT dbg_0i_78_75 (.A(dbg_0_n_78_67),.ZN(dbg_0_dbg_dout[7]));
	NAND2_X1_LVT dbg_0i_78_60 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[6]),.ZN(dbg_0_n_78_54));
	AOI22_X1_LVT dbg_0i_68_13 (.A1(dbg_0_n_68_0),.A2(dbg_mem_din[6]),.B1(dbg_0_n_117),.B2(dbg_mem_din[14]),.ZN(dbg_0_n_68_7));
	INV_X1_LVT dbg_0i_68_14 (.A(dbg_0_n_68_7),.ZN(dbg_0_n_124));
	AOI222_X1_LVT dbg_0i_71_12 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[6]),.B1(dbg_0_n_136),.B2(dbg_reg_din[6]),.C1(dbg_0_n_135),.C2(dbg_0_n_124),.ZN(dbg_0_n_71_6));
	INV_X1_LVT dbg_0i_71_13 (.A(dbg_0_n_71_6),.ZN(dbg_0_n_143));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b6___05F05d (.D(dbg_0_n_143),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[6]),.QN());
	NAND2_X1_LVT dbg_0i_78_61 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[6]),.ZN(dbg_0_n_78_55));
	NAND2_X1_LVT dbg_0i_49_9 (.A1(dbg_0_n_49_4),.A2(dbg_0_n_49_6),.ZN(dbg_0_n_49_9));
	NOR2_X1_LVT dbg_0i_49_24 (.A1(dbg_0_n_49_9),.A2(dbg_0_n_49_20),.ZN(dbg_0_n_93));
	NAND2_X1_LVT dbg_0i_78_62 (.A1(dbg_0_n_93),.A2(dbg_cpu_reset),.ZN(dbg_0_n_78_56));
	NAND2_X1_LVT dbg_0i_78_63 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_57));
	AND4_X1_LVT dbg_0i_78_64 (.A1(dbg_0_n_78_54),.A2(dbg_0_n_78_55),.A3(dbg_0_n_78_56),.A4(dbg_0_n_78_57),.ZN(dbg_0_n_78_58));
	NAND2_X1_LVT dbg_0i_78_65 (.A1(dbg_0_n_91),.A2(cpu_id[6]),.ZN(dbg_0_n_78_59));
	NAND2_X1_LVT dbg_0i_78_66 (.A1(dbg_0_n_99),.A2(1'b0),.ZN(dbg_0_n_78_60));
	NAND2_X1_LVT dbg_0i_78_67 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[6]),.ZN(dbg_0_n_78_61));
	NAND4_X1_LVT dbg_0i_78_68 (.A1(dbg_0_n_78_58),.A2(dbg_0_n_78_59),.A3(dbg_0_n_78_60),.A4(dbg_0_n_78_61),.ZN(dbg_0_dbg_dout[6]));
	NAND2_X1_LVT dbg_0i_78_51 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[5]),.ZN(dbg_0_n_78_46));
	AOI22_X1_LVT dbg_0i_68_11 (.A1(dbg_0_n_68_0),.A2(dbg_mem_din[5]),.B1(dbg_0_n_117),.B2(dbg_mem_din[13]),.ZN(dbg_0_n_68_6));
	INV_X1_LVT dbg_0i_68_12 (.A(dbg_0_n_68_6),.ZN(dbg_0_n_123));
	AOI222_X1_LVT dbg_0i_71_10 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[5]),.B1(dbg_0_n_136),.B2(dbg_reg_din[5]),.C1(dbg_0_n_135),.C2(dbg_0_n_123),.ZN(dbg_0_n_71_5));
	INV_X1_LVT dbg_0i_71_11 (.A(dbg_0_n_71_5),.ZN(dbg_0_n_142));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b5___05F05d (.D(dbg_0_n_142),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[5]),.QN());
	NAND2_X1_LVT dbg_0i_78_52 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[5]),.ZN(dbg_0_n_78_47));
	AND2_X1_LVT dbg_0i_50_0 (.A1(dbg_0_dbg_wr),.A2(dbg_0_n_93),.ZN(dbg_0_cpu_ctl_wr));
	CLKGATETST_X1_LVT dbg_0clk_gate_cpu_ctl_reg___05F_05F0 (.CK(dbg_clk),.E(dbg_0_cpu_ctl_wr),.SE(1'b0),.GCK(dbg_0_n_105));
	DFFS_X1_LVT dbg_0cpu_ctl_reg___05F05b5___05F05d (.D(dbg_0_dbg_din[5]),.SN(dbg_0_n_104),.CK(dbg_0_n_105),.Q(dbg_0_cpu_ctl[2]),.QN());
	NAND2_X1_LVT dbg_0i_78_53 (.A1(dbg_0_n_93),.A2(dbg_0_cpu_ctl[2]),.ZN(dbg_0_n_78_48));
	NAND2_X1_LVT dbg_0i_78_54 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_49));
	AND4_X1_LVT dbg_0i_78_55 (.A1(dbg_0_n_78_46),.A2(dbg_0_n_78_47),.A3(dbg_0_n_78_48),.A4(dbg_0_n_78_49),.ZN(dbg_0_n_78_50));
	NAND2_X1_LVT dbg_0i_78_56 (.A1(dbg_0_n_91),.A2(cpu_id[5]),.ZN(dbg_0_n_78_51));
	NAND2_X1_LVT dbg_0i_78_57 (.A1(dbg_0_n_99),.A2(1'b0),.ZN(dbg_0_n_78_52));
	NAND2_X1_LVT dbg_0i_78_58 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[5]),.ZN(dbg_0_n_78_53));
	NAND4_X1_LVT dbg_0i_78_59 (.A1(dbg_0_n_78_50),.A2(dbg_0_n_78_51),.A3(dbg_0_n_78_52),.A4(dbg_0_n_78_53),.ZN(dbg_0_dbg_dout[5]));
	NAND2_X1_LVT dbg_0i_78_42 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[4]),.ZN(dbg_0_n_78_38));
	AOI22_X1_LVT dbg_0i_68_9 (.A1(dbg_0_n_68_0),.A2(dbg_mem_din[4]),.B1(dbg_0_n_117),.B2(dbg_mem_din[12]),.ZN(dbg_0_n_68_5));
	INV_X1_LVT dbg_0i_68_10 (.A(dbg_0_n_68_5),.ZN(dbg_0_n_122));
	AOI222_X1_LVT dbg_0i_71_8 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[4]),.B1(dbg_0_n_136),.B2(dbg_reg_din[4]),.C1(dbg_0_n_135),.C2(dbg_0_n_122),.ZN(dbg_0_n_71_4));
	INV_X1_LVT dbg_0i_71_9 (.A(dbg_0_n_71_4),.ZN(dbg_0_n_141));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b4___05F05d (.D(dbg_0_n_141),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[4]),.QN());
	NAND2_X1_LVT dbg_0i_78_43 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[4]),.ZN(dbg_0_n_78_39));
	CLKGATETST_X1_LVT dbg_0clk_gate_cpu_ctl_reg___05F_05F1 (.CK(dbg_clk),.E(dbg_0_cpu_ctl_wr),.SE(1'b0),.GCK(dbg_0_n_106));
	DFFS_X1_LVT dbg_0cpu_ctl_reg___05F05b4___05F05d (.D(dbg_0_dbg_din[4]),.SN(dbg_0_n_104),.CK(dbg_0_n_106),.Q(dbg_0_cpu_ctl[1]),.QN());
	NAND2_X1_LVT dbg_0i_78_44 (.A1(dbg_0_n_93),.A2(dbg_0_cpu_ctl[1]),.ZN(dbg_0_n_78_40));
	NAND2_X1_LVT dbg_0i_78_45 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_41));
	AND4_X1_LVT dbg_0i_78_46 (.A1(dbg_0_n_78_38),.A2(dbg_0_n_78_39),.A3(dbg_0_n_78_40),.A4(dbg_0_n_78_41),.ZN(dbg_0_n_78_42));
	NAND2_X1_LVT dbg_0i_78_47 (.A1(dbg_0_n_91),.A2(cpu_id[4]),.ZN(dbg_0_n_78_43));
	NAND2_X1_LVT dbg_0i_78_48 (.A1(dbg_0_n_99),.A2(1'b0),.ZN(dbg_0_n_78_44));
	NAND2_X1_LVT dbg_0i_78_49 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[4]),.ZN(dbg_0_n_78_45));
	NAND4_X1_LVT dbg_0i_78_50 (.A1(dbg_0_n_78_42),.A2(dbg_0_n_78_43),.A3(dbg_0_n_78_44),.A4(dbg_0_n_78_45),.ZN(dbg_0_dbg_dout[4]));
	NAND2_X1_LVT dbg_0i_78_29 (.A1(dbg_0_n_99),.A2(1'b0),.ZN(dbg_0_n_78_26));
	NAND2_X1_LVT dbg_0i_78_30 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[3]),.ZN(dbg_0_n_78_27));
	NAND2_X1_LVT dbg_0i_78_31 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[3]),.ZN(dbg_0_n_78_28));
	AOI22_X1_LVT dbg_0i_68_7 (.A1(dbg_0_n_68_0),.A2(dbg_mem_din[3]),.B1(dbg_0_n_117),.B2(dbg_mem_din[11]),.ZN(dbg_0_n_68_4));
	INV_X1_LVT dbg_0i_68_8 (.A(dbg_0_n_68_4),.ZN(dbg_0_n_121));
	AOI222_X1_LVT dbg_0i_71_6 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[3]),.B1(dbg_0_n_136),.B2(dbg_reg_din[3]),.C1(dbg_0_n_135),.C2(dbg_0_n_121),.ZN(dbg_0_n_71_3));
	INV_X1_LVT dbg_0i_71_7 (.A(dbg_0_n_71_3),.ZN(dbg_0_n_140));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b3___05F05d (.D(dbg_0_n_140),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[3]),.QN());
	NAND2_X1_LVT dbg_0i_78_32 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[3]),.ZN(dbg_0_n_78_29));
	NAND4_X1_LVT dbg_0i_78_33 (.A1(dbg_0_n_78_26),.A2(dbg_0_n_78_27),.A3(dbg_0_n_78_28),.A4(dbg_0_n_78_29),.ZN(dbg_0_n_78_30));
	NAND2_X1_LVT dbg_0i_78_34 (.A1(dbg_0_n_95),.A2(dbg_0_mem_ctl[2]),.ZN(dbg_0_n_78_31));
	NAND2_X1_LVT dbg_0i_49_10 (.A1(dbg_0_n_49_5),.A2(dbg_0_n_49_6),.ZN(dbg_0_n_49_10));
	NOR2_X1_LVT dbg_0i_49_25 (.A1(dbg_0_n_49_10),.A2(dbg_0_n_49_20),.ZN(dbg_0_n_94));
	NAND4_X1_LVT dbg_0i_54_0 (.A1(fe_mdb_in[0]),.A2(fe_mdb_in[1]),.A3(fe_mdb_in[6]),.A4(fe_mdb_in[8]),.ZN(dbg_0_n_54_0));
	CLKGATETST_X1_LVT dbg_0clk_gate_cpu_ctl_reg___05F_05F2 (.CK(dbg_clk),.E(dbg_0_cpu_ctl_wr),.SE(1'b0),.GCK(dbg_0_n_107));
	DFFR_X1_LVT dbg_0cpu_ctl_reg___05F05b3___05F05d (.D(dbg_0_dbg_din[3]),.RN(dbg_0_n_104),.CK(dbg_0_n_107),.Q(dbg_0_cpu_ctl[0]),.QN());
	NAND4_X1_LVT dbg_0i_54_1 (.A1(fe_mdb_in[9]),.A2(fe_mdb_in[14]),.A3(dbg_0_cpu_ctl[0]),.A4(decode_noirq),.ZN(dbg_0_n_54_1));
	NOR4_X1_LVT dbg_0i_54_2 (.A1(dbg_0_n_54_0),.A2(dbg_0_n_54_1),.A3(fe_mdb_in[13]),.A4(fe_mdb_in[15]),.ZN(dbg_0_n_54_2));
	NOR4_X1_LVT dbg_0i_54_3 (.A1(fe_mdb_in[2]),.A2(fe_mdb_in[3]),.A3(fe_mdb_in[4]),.A4(fe_mdb_in[5]),.ZN(dbg_0_n_54_3));
	NOR4_X1_LVT dbg_0i_54_4 (.A1(fe_mdb_in[7]),.A2(fe_mdb_in[10]),.A3(fe_mdb_in[11]),.A4(fe_mdb_in[12]),.ZN(dbg_0_n_54_4));
	AND3_X1_LVT dbg_0i_54_5 (.A1(dbg_0_n_54_2),.A2(dbg_0_n_54_3),.A3(dbg_0_n_54_4),.ZN(dbg_0_dbg_swbrk));
	INV_X1_LVT dbg_0i_76_5 (.A(dbg_0_dbg_din[3]),.ZN(dbg_0_n_76_4));
	AOI21_X1_LVT dbg_0i_76_6 (.A(dbg_0_dbg_swbrk),.B1(dbg_0_n_76_4),.B2(dbg_0_cpu_stat[1]),.ZN(dbg_0_n_76_5));
	AND2_X1_LVT dbg_0i_50_1 (.A1(dbg_0_dbg_wr),.A2(dbg_0_n_94),.ZN(dbg_0_n_100));
	INV_X1_LVT dbg_0i_76_2 (.A(dbg_0_n_100),.ZN(dbg_0_n_76_2));
	NOR2_X1_LVT dbg_0i_76_7 (.A1(dbg_0_cpu_stat[1]),.A2(dbg_0_dbg_swbrk),.ZN(dbg_0_n_76_6));
	OAI22_X1_LVT dbg_0i_76_8 (.A1(dbg_0_n_76_5),.A2(dbg_0_n_76_2),.B1(dbg_0_n_76_6),.B2(dbg_0_n_100),.ZN(dbg_0_n_155));
	DFFR_X1_LVT dbg_0cpu_stat_reg___05F05b3___05F05d (.D(dbg_0_n_155),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_cpu_stat[1]),.QN());
	NAND2_X1_LVT dbg_0i_78_35 (.A1(dbg_0_n_94),.A2(dbg_0_cpu_stat[1]),.ZN(dbg_0_n_78_32));
	NAND2_X1_LVT dbg_0i_78_36 (.A1(dbg_0_n_93),.A2(dbg_0_cpu_ctl[0]),.ZN(dbg_0_n_78_33));
	NAND2_X1_LVT dbg_0i_78_37 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_34));
	NAND4_X1_LVT dbg_0i_78_38 (.A1(dbg_0_n_78_31),.A2(dbg_0_n_78_32),.A3(dbg_0_n_78_33),.A4(dbg_0_n_78_34),.ZN(dbg_0_n_78_35));
	NOR2_X1_LVT dbg_0i_78_39 (.A1(dbg_0_n_78_30),.A2(dbg_0_n_78_35),.ZN(dbg_0_n_78_36));
	NAND2_X1_LVT dbg_0i_78_40 (.A1(dbg_0_n_91),.A2(cpu_id[3]),.ZN(dbg_0_n_78_37));
	NAND2_X1_LVT dbg_0i_78_41 (.A1(dbg_0_n_78_36),.A2(dbg_0_n_78_37),.ZN(dbg_0_dbg_dout[3]));
	NAND2_X1_LVT dbg_0i_78_18 (.A1(dbg_0_n_91),.A2(cpu_id[2]),.ZN(dbg_0_n_78_16));
	NAND2_X1_LVT dbg_0i_78_19 (.A1(dbg_0_n_99),.A2(1'b0),.ZN(dbg_0_n_78_17));
	NAND2_X1_LVT dbg_0i_78_20 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[2]),.ZN(dbg_0_n_78_18));
	NAND2_X1_LVT dbg_0i_78_21 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[2]),.ZN(dbg_0_n_78_19));
	NAND4_X1_LVT dbg_0i_78_22 (.A1(dbg_0_n_78_16),.A2(dbg_0_n_78_17),.A3(dbg_0_n_78_18),.A4(dbg_0_n_78_19),.ZN(dbg_0_n_78_20));
	AOI22_X1_LVT dbg_0i_68_5 (.A1(dbg_0_n_68_0),.A2(dbg_mem_din[2]),.B1(dbg_0_n_117),.B2(dbg_mem_din[10]),.ZN(dbg_0_n_68_3));
	INV_X1_LVT dbg_0i_68_6 (.A(dbg_0_n_68_3),.ZN(dbg_0_n_120));
	AOI222_X1_LVT dbg_0i_71_4 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[2]),.B1(dbg_0_n_136),.B2(dbg_reg_din[2]),.C1(dbg_0_n_135),.C2(dbg_0_n_120),.ZN(dbg_0_n_71_2));
	INV_X1_LVT dbg_0i_71_5 (.A(dbg_0_n_71_2),.ZN(dbg_0_n_139));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b2___05F05d (.D(dbg_0_n_139),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[2]),.QN());
	NAND2_X1_LVT dbg_0i_78_23 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[2]),.ZN(dbg_0_n_78_21));
	NAND2_X1_LVT dbg_0i_78_24 (.A1(dbg_0_n_95),.A2(dbg_0_mem_ctl[1]),.ZN(dbg_0_n_78_22));
	INV_X1_LVT dbg_0i_76_0 (.A(dbg_0_dbg_din[2]),.ZN(dbg_0_n_76_0));
	AOI21_X1_LVT dbg_0i_76_1 (.A(puc_pnd_set),.B1(dbg_0_n_76_0),.B2(dbg_0_cpu_stat[0]),.ZN(dbg_0_n_76_1));
	NOR2_X1_LVT dbg_0i_76_3 (.A1(dbg_0_cpu_stat[0]),.A2(puc_pnd_set),.ZN(dbg_0_n_76_3));
	OAI22_X1_LVT dbg_0i_76_4 (.A1(dbg_0_n_76_1),.A2(dbg_0_n_76_2),.B1(dbg_0_n_76_3),.B2(dbg_0_n_100),.ZN(dbg_0_n_154));
	DFFR_X1_LVT dbg_0cpu_stat_reg___05F05b2___05F05d (.D(dbg_0_n_154),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_cpu_stat[0]),.QN());
	NAND2_X1_LVT dbg_0i_78_25 (.A1(dbg_0_n_94),.A2(dbg_0_cpu_stat[0]),.ZN(dbg_0_n_78_23));
	NAND2_X1_LVT dbg_0i_78_26 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_24));
	NAND4_X1_LVT dbg_0i_78_27 (.A1(dbg_0_n_78_21),.A2(dbg_0_n_78_22),.A3(dbg_0_n_78_23),.A4(dbg_0_n_78_24),.ZN(dbg_0_n_78_25));
	OR2_X1_LVT dbg_0i_78_28 (.A1(dbg_0_n_78_20),.A2(dbg_0_n_78_25),.ZN(dbg_0_dbg_dout[2]));
	NAND2_X1_LVT dbg_0i_78_9 (.A1(dbg_0_n_96),.A2(dbg_mem_addr[1]),.ZN(dbg_0_n_78_8));
	AOI22_X1_LVT dbg_0i_68_3 (.A1(dbg_0_n_68_0),.A2(dbg_mem_din[1]),.B1(dbg_0_n_117),.B2(dbg_mem_din[9]),.ZN(dbg_0_n_68_2));
	INV_X1_LVT dbg_0i_68_4 (.A(dbg_0_n_68_2),.ZN(dbg_0_n_119));
	AOI222_X1_LVT dbg_0i_71_2 (.A1(dbg_0_mem_data_wr),.A2(dbg_0_dbg_din[1]),.B1(dbg_0_n_136),.B2(dbg_reg_din[1]),.C1(dbg_0_n_135),.C2(dbg_0_n_119),.ZN(dbg_0_n_71_1));
	INV_X1_LVT dbg_0i_71_3 (.A(dbg_0_n_71_1),.ZN(dbg_0_n_138));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b1___05F05d (.D(dbg_0_n_138),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[1]),.QN());
	NAND2_X1_LVT dbg_0i_78_10 (.A1(dbg_0_n_97),.A2(dbg_0_mem_data[1]),.ZN(dbg_0_n_78_9));
	NAND2_X1_LVT dbg_0i_78_11 (.A1(dbg_0_n_95),.A2(dbg_0_mem_ctl[0]),.ZN(dbg_0_n_78_10));
	NAND2_X1_LVT dbg_0i_78_12 (.A1(dbg_0_n_92),.A2(cpu_id[0]),.ZN(dbg_0_n_78_11));
	AND4_X1_LVT dbg_0i_78_13 (.A1(dbg_0_n_78_8),.A2(dbg_0_n_78_9),.A3(dbg_0_n_78_10),.A4(dbg_0_n_78_11),.ZN(dbg_0_n_78_12));
	NAND2_X1_LVT dbg_0i_78_14 (.A1(dbg_0_n_91),.A2(cpu_id[1]),.ZN(dbg_0_n_78_13));
	NAND2_X1_LVT dbg_0i_78_15 (.A1(dbg_0_n_99),.A2(1'b0),.ZN(dbg_0_n_78_14));
	NAND2_X1_LVT dbg_0i_78_16 (.A1(dbg_0_n_98),.A2(dbg_0_mem_cnt[1]),.ZN(dbg_0_n_78_15));
	NAND4_X1_LVT dbg_0i_78_17 (.A1(dbg_0_n_78_12),.A2(dbg_0_n_78_13),.A3(dbg_0_n_78_14),.A4(dbg_0_n_78_15),.ZN(dbg_0_dbg_dout[1]));
	NAND2_X1_LVT dbg_0i_78_0 (.A1(dbg_mem_addr[0]),.A2(dbg_0_n_96),.ZN(dbg_0_n_78_0));
	AOI22_X1_LVT dbg_0i_68_1 (.A1(dbg_0_n_68_0),.A2(dbg_mem_din[0]),.B1(dbg_mem_din[8]),.B2(dbg_0_n_117),.ZN(dbg_0_n_68_1));
	INV_X1_LVT dbg_0i_68_2 (.A(dbg_0_n_68_1),.ZN(dbg_0_n_118));
	AOI222_X1_LVT dbg_0i_71_0 (.A1(dbg_0_dbg_din[0]),.A2(dbg_0_mem_data_wr),.B1(dbg_reg_din[0]),.B2(dbg_0_n_136),.C1(dbg_0_n_118),.C2(dbg_0_n_135),.ZN(dbg_0_n_71_0));
	INV_X1_LVT dbg_0i_71_1 (.A(dbg_0_n_71_0),.ZN(dbg_0_n_137));
	DFFR_X1_LVT dbg_0mem_data_reg___05F05b0___05F05d (.D(dbg_0_n_137),.RN(dbg_0_n_104),.CK(dbg_0_n_134),.Q(dbg_0_mem_data[0]),.QN());
	NAND2_X1_LVT dbg_0i_78_1 (.A1(dbg_0_mem_data[0]),.A2(dbg_0_n_97),.ZN(dbg_0_n_78_1));
	NAND2_X1_LVT dbg_0i_78_2 (.A1(cpu_halt_st),.A2(dbg_0_n_94),.ZN(dbg_0_n_78_2));
	NAND2_X1_LVT dbg_0i_78_3 (.A1(cpu_id[0]),.A2(dbg_0_n_92),.ZN(dbg_0_n_78_3));
	AND4_X1_LVT dbg_0i_78_4 (.A1(dbg_0_n_78_0),.A2(dbg_0_n_78_1),.A3(dbg_0_n_78_2),.A4(dbg_0_n_78_3),.ZN(dbg_0_n_78_4));
	NAND2_X1_LVT dbg_0i_78_5 (.A1(cpu_id[0]),.A2(dbg_0_n_91),.ZN(dbg_0_n_78_5));
	NAND2_X1_LVT dbg_0i_78_6 (.A1(1'b0),.A2(dbg_0_n_99),.ZN(dbg_0_n_78_6));
	NAND2_X1_LVT dbg_0i_78_7 (.A1(dbg_0_mem_cnt[0]),.A2(dbg_0_n_98),.ZN(dbg_0_n_78_7));
	NAND4_X1_LVT dbg_0i_78_8 (.A1(dbg_0_n_78_4),.A2(dbg_0_n_78_5),.A3(dbg_0_n_78_6),.A4(dbg_0_n_78_7),.ZN(dbg_0_dbg_dout[0]));
	AND2_X1_LVT dbg_0i_79_0 (.A1(dbg_0_mem_ctl[0]),.A2(dbg_0_mem_burst_start),.ZN(dbg_0_mem_burst_wr));
	INV_X1_LVT dbg_0dbg_uart_0i_4_0 (.A(dbg_0_dbg_rd_rdy),.ZN(dbg_0_dbg_uart_0_n_4_0));
	INV_X1_LVT dbg_0dbg_uart_0i_57_0 (.A(dbg_uart_rxd),.ZN(dbg_0_dbg_uart_0_n_136));
	INV_X1_LVT dbg_0dbg_uart_0sync_cell_uart_rxdi_0_0 (.A(dbg_rst),.ZN(dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_0));
	DFFR_X1_LVT dbg_0dbg_uart_0sync_cell_uart_rxddata_sync_reg___05F05b0___05F05d (.D(dbg_0_dbg_uart_0_n_136),.RN(dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_0),.CK(dbg_clk),.Q(dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_1),.QN());
	DFFR_X1_LVT dbg_0dbg_uart_0sync_cell_uart_rxddata_sync_reg___05F05b1___05F05d (.D(dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_1),.RN(dbg_0_dbg_uart_0_sync_cell_uart_rxd_n_0),.CK(dbg_clk),.Q(dbg_0_dbg_uart_0_uart_rxd_n),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_0_0 (.A(dbg_0_dbg_uart_0_uart_rxd_n),.ZN(dbg_0_dbg_uart_0_uart_rxd));
	INV_X1_LVT dbg_0dbg_uart_0i_2_0 (.A(dbg_0_dbg_uart_0_uart_rxd),.ZN(dbg_0_dbg_uart_0_n_2_0));
	INV_X1_LVT dbg_0dbg_uart_0i_46_0 (.A(dbg_rst),.ZN(dbg_0_dbg_uart_0_n_130));
	DFFS_X1_LVT dbg_0dbg_uart_0rxd_buf_reg___05F05b0___05F05d (.D(dbg_0_dbg_uart_0_uart_rxd),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_clk),.Q(dbg_0_dbg_uart_0_rxd_buf[0]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_2_1 (.A(dbg_0_dbg_uart_0_rxd_buf[0]),.ZN(dbg_0_dbg_uart_0_n_2_1));
	DFFS_X1_LVT dbg_0dbg_uart_0rxd_buf_reg___05F05b1___05F05d (.D(dbg_0_dbg_uart_0_rxd_buf[0]),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_clk),.Q(dbg_0_dbg_uart_0_rxd_buf[1]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_2_2 (.A(dbg_0_dbg_uart_0_rxd_buf[1]),.ZN(dbg_0_dbg_uart_0_n_2_2));
	OAI222_X1_LVT dbg_0dbg_uart_0i_2_3 (.A1(dbg_0_dbg_uart_0_n_2_0),.A2(dbg_0_dbg_uart_0_n_2_1),.B1(dbg_0_dbg_uart_0_n_2_1),.B2(dbg_0_dbg_uart_0_n_2_2),.C1(dbg_0_dbg_uart_0_n_2_0),.C2(dbg_0_dbg_uart_0_n_2_2),.ZN(dbg_0_dbg_uart_0_rxd_maj_nxt));
	DFFS_X1_LVT dbg_0dbg_uart_0rxd_maj_reg (.D(dbg_0_dbg_uart_0_rxd_maj_nxt),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_clk),.Q(dbg_0_dbg_uart_0_rxd_maj),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_4_36 (.A(dbg_0_dbg_uart_0_rxd_maj),.ZN(dbg_0_dbg_uart_0_n_4_18));
	NAND2_X1_LVT dbg_0dbg_uart_0i_4_37 (.A1(dbg_0_dbg_uart_0_n_4_18),.A2(dbg_0_dbg_uart_0_n_4_0),.ZN(dbg_0_dbg_uart_0_n_19));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F16 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_53));
	DFFR_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b1___05F05d (.D(dbg_0_dbg_uart_0_n_58),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_53),.Q(dbg_0_dbg_uart_0_n_54),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_21_0 (.A(dbg_0_dbg_uart_0_n_56),.ZN(dbg_0_dbg_uart_0_n_57));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F17 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_55));
	DFFR_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b0___05F05d (.D(dbg_0_dbg_uart_0_n_57),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_55),.Q(dbg_0_dbg_uart_0_n_56),.QN());
	HA_X1_LVT dbg_0dbg_uart_0i_21_1 (.A(dbg_0_dbg_uart_0_n_54),.B(dbg_0_dbg_uart_0_n_56),.CO(dbg_0_dbg_uart_0_n_21_0),.S(dbg_0_dbg_uart_0_n_58));
	HA_X1_LVT dbg_0dbg_uart_0i_21_2 (.A(dbg_0_dbg_uart_0_n_52),.B(dbg_0_dbg_uart_0_n_21_0),.CO(dbg_0_dbg_uart_0_n_21_1),.S(dbg_0_dbg_uart_0_n_59));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F15 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_51));
	DFFR_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b2___05F05d (.D(dbg_0_dbg_uart_0_n_59),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_51),.Q(dbg_0_dbg_uart_0_n_52),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_22_1 (.A(dbg_0_dbg_uart_0_n_52),.ZN(dbg_0_dbg_uart_0_n_22_1));
	NOR3_X1_LVT dbg_0dbg_uart_0i_8_4 (.A1(dbg_0_dbg_uart_0_n_8_3),.A2(dbg_0_dbg_uart_0_uart_state[0]),.A3(dbg_0_dbg_uart_0_uart_state[1]),.ZN(dbg_0_dbg_uart_0_n_8_4));
	INV_X1_LVT dbg_0dbg_uart_0i_8_5 (.A(dbg_0_dbg_uart_0_n_8_4),.ZN(dbg_0_dbg_uart_0_n_8_5));
	NAND3_X1_LVT dbg_0dbg_uart_0i_8_7 (.A1(dbg_0_dbg_uart_0_n_8_0),.A2(dbg_0_dbg_uart_0_uart_state[0]),.A3(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_8_7));
	INV_X1_LVT dbg_0dbg_uart_0i_7_0 (.A(dbg_0_mem_burst),.ZN(dbg_0_dbg_uart_0_n_7_0));
	NOR2_X1_LVT dbg_0dbg_uart_0i_7_1 (.A1(dbg_0_dbg_uart_0_n_7_0),.A2(dbg_0_mem_burst_end),.ZN(dbg_0_dbg_uart_0_n_22));
	INV_X1_LVT dbg_0dbg_uart_0i_8_27 (.A(dbg_0_dbg_uart_0_n_22),.ZN(dbg_0_dbg_uart_0_n_8_26));
	INV_X1_LVT dbg_0dbg_uart_0i_8_20 (.A(dbg_0_mem_burst_wr),.ZN(dbg_0_dbg_uart_0_n_8_20));
	NAND2_X1_LVT dbg_0dbg_uart_0i_8_21 (.A1(dbg_0_dbg_uart_0_n_8_20),.A2(dbg_0_mem_burst_rd),.ZN(dbg_0_dbg_uart_0_n_8_21));
	INV_X1_LVT dbg_0dbg_uart_0i_8_29 (.A(dbg_0_dbg_uart_0_n_8_21),.ZN(dbg_0_dbg_uart_0_n_8_27));
	OR2_X1_LVT dbg_0dbg_uart_0i_8_15 (.A1(dbg_0_mem_burst_rd),.A2(dbg_0_mem_burst_wr),.ZN(dbg_0_dbg_uart_0_n_8_15));
	NOR2_X1_LVT dbg_0dbg_uart_0i_8_16 (.A1(dbg_0_dbg_uart_0_n_8_15),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.ZN(dbg_0_dbg_uart_0_n_8_16));
	AND2_X1_LVT dbg_0dbg_uart_0i_8_17 (.A1(dbg_0_dbg_uart_0_n_8_16),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.ZN(dbg_0_dbg_uart_0_n_8_17));
	INV_X1_LVT dbg_0dbg_uart_0i_8_30 (.A(dbg_0_dbg_uart_0_xfer_buf[0]),.ZN(dbg_0_dbg_uart_0_n_8_28));
	AOI211_X1_LVT dbg_0dbg_uart_0i_8_31 (.A(dbg_0_dbg_uart_0_n_8_27),.B(dbg_0_dbg_uart_0_n_8_17),.C1(dbg_0_dbg_uart_0_n_8_16),.C2(dbg_0_dbg_uart_0_n_8_28),.ZN(dbg_0_dbg_uart_0_n_8_29));
	INV_X1_LVT dbg_0dbg_uart_0i_8_24 (.A(dbg_0_dbg_uart_0_n_8_10),.ZN(dbg_0_dbg_uart_0_n_8_24));
	OAI221_X1_LVT dbg_0dbg_uart_0i_8_32 (.A(dbg_0_dbg_uart_0_n_8_5),.B1(dbg_0_dbg_uart_0_n_8_7),.B2(dbg_0_dbg_uart_0_n_8_26),.C1(dbg_0_dbg_uart_0_n_8_29),.C2(dbg_0_dbg_uart_0_n_8_24),.ZN(dbg_0_dbg_uart_0_uart_state_nxt_reg[2]));
	INV_X1_LVT dbg_0dbg_uart_0i_39_0 (.A(dbg_0_dbg_uart_0_xfer_bit[0]),.ZN(dbg_0_dbg_uart_0_n_119));
	AOI21_X1_LVT dbg_0dbg_uart_0i_41_1 (.A(dbg_0_dbg_uart_0_n_123),.B1(dbg_0_dbg_uart_0_n_41_0),.B2(dbg_0_dbg_uart_0_n_119),.ZN(dbg_0_dbg_uart_0_n_41_1));
	INV_X1_LVT dbg_0dbg_uart_0i_41_2 (.A(dbg_0_dbg_uart_0_n_41_1),.ZN(dbg_0_dbg_uart_0_n_124));
	INV_X1_LVT dbg_0dbg_uart_0i_42_0 (.A(dbg_0_dbg_uart_0_xfer_done),.ZN(dbg_0_dbg_uart_0_n_42_0));
	INV_X1_LVT dbg_0dbg_uart_0i_42_1 (.A(dbg_0_dbg_uart_0_n_123),.ZN(dbg_0_dbg_uart_0_n_42_1));
	NAND3_X1_LVT dbg_0dbg_uart_0i_42_2 (.A1(dbg_0_dbg_uart_0_n_42_0),.A2(dbg_0_dbg_uart_0_n_42_1),.A3(dbg_0_dbg_uart_0_xfer_bit_inc),.ZN(dbg_0_dbg_uart_0_n_42_2));
	NAND3_X1_LVT dbg_0dbg_uart_0i_42_3 (.A1(dbg_0_dbg_uart_0_n_42_2),.A2(dbg_0_dbg_uart_0_n_42_0),.A3(dbg_0_dbg_uart_0_n_42_1),.ZN(dbg_0_dbg_uart_0_n_128));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_xfer_bit_reg (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_128),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_118));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_bit_reg___05F05b0___05F05d (.D(dbg_0_dbg_uart_0_n_124),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_118),.Q(dbg_0_dbg_uart_0_xfer_bit[0]),.QN());
	HA_X1_LVT dbg_0dbg_uart_0i_39_1 (.A(dbg_0_dbg_uart_0_xfer_bit[1]),.B(dbg_0_dbg_uart_0_xfer_bit[0]),.CO(dbg_0_dbg_uart_0_n_39_0),.S(dbg_0_dbg_uart_0_n_120));
	AND2_X1_LVT dbg_0dbg_uart_0i_41_3 (.A1(dbg_0_dbg_uart_0_n_41_0),.A2(dbg_0_dbg_uart_0_n_120),.ZN(dbg_0_dbg_uart_0_n_125));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_bit_reg___05F05b1___05F05d (.D(dbg_0_dbg_uart_0_n_125),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_118),.Q(dbg_0_dbg_uart_0_xfer_bit[1]),.QN());
	HA_X1_LVT dbg_0dbg_uart_0i_39_2 (.A(dbg_0_dbg_uart_0_xfer_bit[2]),.B(dbg_0_dbg_uart_0_n_39_0),.CO(dbg_0_dbg_uart_0_n_39_1),.S(dbg_0_dbg_uart_0_n_121));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_39_3 (.A(dbg_0_dbg_uart_0_xfer_bit[3]),.B(dbg_0_dbg_uart_0_n_39_1),.ZN(dbg_0_dbg_uart_0_n_39_2));
	INV_X1_LVT dbg_0dbg_uart_0i_39_4 (.A(dbg_0_dbg_uart_0_n_39_2),.ZN(dbg_0_dbg_uart_0_n_122));
	AND2_X1_LVT dbg_0dbg_uart_0i_41_5 (.A1(dbg_0_dbg_uart_0_n_41_0),.A2(dbg_0_dbg_uart_0_n_122),.ZN(dbg_0_dbg_uart_0_n_127));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_bit_reg___05F05b3___05F05d (.D(dbg_0_dbg_uart_0_n_127),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_118),.Q(dbg_0_dbg_uart_0_xfer_bit[3]),.QN());
	NOR4_X1_LVT dbg_0dbg_uart_0i_36_0 (.A1(dbg_0_dbg_uart_0_xfer_bit[0]),.A2(dbg_0_dbg_uart_0_xfer_bit[1]),.A3(dbg_0_dbg_uart_0_xfer_bit[2]),.A4(dbg_0_dbg_uart_0_xfer_bit[3]),.ZN(dbg_0_dbg_uart_0_n_116));
	OR3_X1_LVT dbg_0dbg_uart_0i_37_0 (.A1(dbg_0_dbg_uart_0_uart_state[0]),.A2(dbg_0_dbg_uart_0_uart_state[1]),.A3(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_117));
	INV_X1_LVT dbg_0dbg_uart_0i_15_0 (.A(dbg_0_dbg_uart_0_rxd_maj),.ZN(dbg_0_dbg_uart_0_n_15_0));
	NOR2_X1_LVT dbg_0dbg_uart_0i_15_1 (.A1(dbg_0_dbg_uart_0_n_15_0),.A2(dbg_0_dbg_uart_0_rxd_maj_nxt),.ZN(dbg_0_dbg_uart_0_rxd_fe));
	AND3_X1_LVT dbg_0dbg_uart_0i_40_0 (.A1(dbg_0_dbg_uart_0_n_116),.A2(dbg_0_dbg_uart_0_n_117),.A3(dbg_0_dbg_uart_0_rxd_fe),.ZN(dbg_0_dbg_uart_0_n_40_0));
	INV_X1_LVT dbg_0dbg_uart_0i_13_5 (.A(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_13_2));
	NOR3_X1_LVT dbg_0dbg_uart_0i_13_6 (.A1(dbg_0_dbg_uart_0_n_13_2),.A2(dbg_0_dbg_uart_0_uart_state[0]),.A3(dbg_0_dbg_uart_0_uart_state[1]),.ZN(dbg_0_dbg_uart_0_n_28));
	AOI21_X1_LVT dbg_0dbg_uart_0i_24_0 (.A(dbg_0_dbg_rd_rdy),.B1(dbg_0_dbg_uart_0_xfer_done),.B2(dbg_0_dbg_uart_0_n_28),.ZN(dbg_0_dbg_uart_0_n_24_0));
	INV_X1_LVT dbg_0dbg_uart_0i_24_1 (.A(dbg_0_dbg_uart_0_n_24_0),.ZN(dbg_0_dbg_uart_0_txd_start));
	OR2_X1_LVT dbg_0dbg_uart_0i_40_1 (.A1(dbg_0_dbg_uart_0_n_40_0),.A2(dbg_0_dbg_uart_0_txd_start),.ZN(dbg_0_dbg_uart_0_n_123));
	NOR2_X1_LVT dbg_0dbg_uart_0i_41_0 (.A1(dbg_0_dbg_uart_0_xfer_done),.A2(dbg_0_dbg_uart_0_n_123),.ZN(dbg_0_dbg_uart_0_n_41_0));
	AND2_X1_LVT dbg_0dbg_uart_0i_41_4 (.A1(dbg_0_dbg_uart_0_n_41_0),.A2(dbg_0_dbg_uart_0_n_121),.ZN(dbg_0_dbg_uart_0_n_126));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_bit_reg___05F05b2___05F05d (.D(dbg_0_dbg_uart_0_n_126),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_118),.Q(dbg_0_dbg_uart_0_xfer_bit[2]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_44_0 (.A(dbg_0_dbg_uart_0_xfer_bit[2]),.ZN(dbg_0_dbg_uart_0_n_44_0));
	INV_X1_LVT dbg_0dbg_uart_0i_13_0 (.A(dbg_0_dbg_uart_0_uart_state[1]),.ZN(dbg_0_dbg_uart_0_n_13_0));
	NOR3_X1_LVT dbg_0dbg_uart_0i_13_1 (.A1(dbg_0_dbg_uart_0_n_13_0),.A2(dbg_0_dbg_uart_0_uart_state[0]),.A3(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_25));
	INV_X1_LVT dbg_0dbg_uart_0i_13_2 (.A(dbg_0_dbg_uart_0_uart_state[0]),.ZN(dbg_0_dbg_uart_0_n_13_1));
	NOR3_X1_LVT dbg_0dbg_uart_0i_13_4 (.A1(dbg_0_dbg_uart_0_n_13_1),.A2(dbg_0_dbg_uart_0_uart_state[1]),.A3(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_27));
	NOR3_X1_LVT dbg_0dbg_uart_0i_13_3 (.A1(dbg_0_dbg_uart_0_n_13_0),.A2(dbg_0_dbg_uart_0_n_13_1),.A3(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_26));
	OR3_X1_LVT dbg_0dbg_uart_0i_25_0 (.A1(dbg_0_dbg_uart_0_n_25),.A2(dbg_0_dbg_uart_0_n_27),.A3(dbg_0_dbg_uart_0_n_26),.ZN(dbg_0_dbg_uart_0_rx_active));
	NAND4_X1_LVT dbg_0dbg_uart_0i_44_1 (.A1(dbg_0_dbg_uart_0_n_44_0),.A2(dbg_0_dbg_uart_0_xfer_bit[1]),.A3(dbg_0_dbg_uart_0_xfer_bit[3]),.A4(dbg_0_dbg_uart_0_rx_active),.ZN(dbg_0_dbg_uart_0_n_44_1));
	INV_X1_LVT dbg_0dbg_uart_0i_44_2 (.A(dbg_0_dbg_uart_0_rx_active),.ZN(dbg_0_dbg_uart_0_n_44_2));
	NAND4_X1_LVT dbg_0dbg_uart_0i_44_3 (.A1(dbg_0_dbg_uart_0_n_44_2),.A2(dbg_0_dbg_uart_0_xfer_bit[0]),.A3(dbg_0_dbg_uart_0_xfer_bit[1]),.A4(dbg_0_dbg_uart_0_xfer_bit[3]),.ZN(dbg_0_dbg_uart_0_n_44_3));
	OAI22_X1_LVT dbg_0dbg_uart_0i_44_4 (.A1(dbg_0_dbg_uart_0_n_44_1),.A2(dbg_0_dbg_uart_0_xfer_bit[0]),.B1(dbg_0_dbg_uart_0_n_44_3),.B2(dbg_0_dbg_uart_0_xfer_bit[2]),.ZN(dbg_0_dbg_uart_0_xfer_done));
	NOR3_X1_LVT dbg_0dbg_uart_0i_11_0 (.A1(dbg_0_dbg_uart_0_xfer_done),.A2(dbg_0_mem_burst_rd),.A3(dbg_0_mem_burst_wr),.ZN(dbg_0_dbg_uart_0_n_11_0));
	NAND2_X1_LVT dbg_0dbg_uart_0i_14_0 (.A1(dbg_0_dbg_uart_0_n_29),.A2(dbg_0_dbg_uart_0_rxd_maj_nxt),.ZN(dbg_0_dbg_uart_0_n_14_0));
	NOR2_X1_LVT dbg_0dbg_uart_0i_14_1 (.A1(dbg_0_dbg_uart_0_n_14_0),.A2(dbg_0_dbg_uart_0_rxd_maj),.ZN(dbg_0_dbg_uart_0_n_31));
	NAND2_X1_LVT dbg_0dbg_uart_0i_11_1 (.A1(dbg_0_dbg_uart_0_n_31),.A2(dbg_0_dbg_uart_0_sync_busy),.ZN(dbg_0_dbg_uart_0_n_11_1));
	NAND2_X1_LVT dbg_0dbg_uart_0i_11_2 (.A1(dbg_0_dbg_uart_0_n_11_0),.A2(dbg_0_dbg_uart_0_n_11_1),.ZN(dbg_0_dbg_uart_0_n_24));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_uart_state_reg (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_24),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_23));
	DFFR_X1_LVT dbg_0dbg_uart_0uart_state_reg___05F05b2___05F05d (.D(dbg_0_dbg_uart_0_uart_state_nxt_reg[2]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_23),.Q(dbg_0_dbg_uart_0_uart_state[2]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_8_3 (.A(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_8_3));
	AND3_X1_LVT dbg_0dbg_uart_0i_8_10 (.A1(dbg_0_dbg_uart_0_n_8_0),.A2(dbg_0_dbg_uart_0_n_8_3),.A3(dbg_0_dbg_uart_0_uart_state[0]),.ZN(dbg_0_dbg_uart_0_n_8_10));
	INV_X1_LVT dbg_0dbg_uart_0i_8_18 (.A(dbg_0_dbg_uart_0_xfer_buf[0]),.ZN(dbg_0_dbg_uart_0_n_8_18));
	NOR2_X1_LVT dbg_0dbg_uart_0i_8_19 (.A1(dbg_0_dbg_uart_0_n_8_15),.A2(dbg_0_dbg_uart_0_n_8_18),.ZN(dbg_0_dbg_uart_0_n_8_19));
	OAI21_X1_LVT dbg_0dbg_uart_0i_8_26 (.A(dbg_0_dbg_uart_0_n_8_10),.B1(dbg_0_dbg_uart_0_n_8_19),.B2(dbg_0_mem_burst_wr),.ZN(dbg_0_dbg_uart_0_n_8_25));
	NAND3_X1_LVT dbg_0dbg_uart_0i_8_6 (.A1(dbg_0_dbg_uart_0_n_8_3),.A2(dbg_0_dbg_uart_0_uart_state[0]),.A3(dbg_0_dbg_uart_0_uart_state[1]),.ZN(dbg_0_dbg_uart_0_n_8_6));
	OAI211_X1_LVT dbg_0dbg_uart_0i_8_28 (.A(dbg_0_dbg_uart_0_n_8_25),.B(dbg_0_dbg_uart_0_n_8_2),.C1(dbg_0_dbg_uart_0_n_8_6),.C2(dbg_0_dbg_uart_0_n_8_26),.ZN(dbg_0_dbg_uart_0_uart_state_nxt_reg[1]));
	DFFR_X1_LVT dbg_0dbg_uart_0uart_state_reg___05F05b1___05F05d (.D(dbg_0_dbg_uart_0_uart_state_nxt_reg[1]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_23),.Q(dbg_0_dbg_uart_0_uart_state[1]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_8_0 (.A(dbg_0_dbg_uart_0_uart_state[1]),.ZN(dbg_0_dbg_uart_0_n_8_0));
	NOR3_X1_LVT dbg_0dbg_uart_0i_8_1 (.A1(dbg_0_dbg_uart_0_n_8_0),.A2(dbg_0_dbg_uart_0_uart_state[0]),.A3(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_8_1));
	INV_X1_LVT dbg_0dbg_uart_0i_8_2 (.A(dbg_0_dbg_uart_0_n_8_1),.ZN(dbg_0_dbg_uart_0_n_8_2));
	NAND4_X1_LVT dbg_0dbg_uart_0i_8_8 (.A1(dbg_0_dbg_uart_0_n_8_2),.A2(dbg_0_dbg_uart_0_n_8_5),.A3(dbg_0_dbg_uart_0_n_8_6),.A4(dbg_0_dbg_uart_0_n_8_7),.ZN(dbg_0_dbg_uart_0_n_8_8));
	NOR3_X1_LVT dbg_0dbg_uart_0i_8_9 (.A1(dbg_0_dbg_uart_0_uart_state[0]),.A2(dbg_0_dbg_uart_0_uart_state[1]),.A3(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_8_9));
	OR3_X1_LVT dbg_0dbg_uart_0i_8_11 (.A1(dbg_0_dbg_uart_0_n_8_8),.A2(dbg_0_dbg_uart_0_n_8_9),.A3(dbg_0_dbg_uart_0_n_8_10),.ZN(dbg_0_dbg_uart_0_n_8_11));
	NAND2_X1_LVT dbg_0dbg_uart_0i_8_12 (.A1(dbg_0_mem_ctl[2]),.A2(dbg_0_dbg_uart_0_n_22),.ZN(dbg_0_dbg_uart_0_n_8_12));
	AOI22_X1_LVT dbg_0dbg_uart_0i_8_13 (.A1(dbg_0_dbg_uart_0_n_8_6),.A2(dbg_0_dbg_uart_0_n_8_7),.B1(dbg_0_dbg_uart_0_n_8_12),.B2(dbg_0_dbg_uart_0_n_22),.ZN(dbg_0_dbg_uart_0_n_8_13));
	NOR4_X1_LVT dbg_0dbg_uart_0i_8_14 (.A1(dbg_0_dbg_uart_0_n_8_13),.A2(dbg_0_dbg_uart_0_n_8_4),.A3(dbg_0_dbg_uart_0_n_8_1),.A4(dbg_0_dbg_uart_0_n_8_9),.ZN(dbg_0_dbg_uart_0_n_8_14));
	NAND2_X1_LVT dbg_0dbg_uart_0i_8_22 (.A1(dbg_0_dbg_uart_0_n_8_21),.A2(dbg_0_dbg_uart_0_n_8_20),.ZN(dbg_0_dbg_uart_0_n_8_22));
	AOI221_X1_LVT dbg_0dbg_uart_0i_8_23 (.A(dbg_0_dbg_uart_0_n_8_17),.B1(dbg_0_dbg_uart_0_n_8_19),.B2(dbg_0_dbg_uart_0_xfer_buf[0]),.C1(dbg_0_dbg_uart_0_n_8_22),.C2(dbg_0_mem_ctl[2]),.ZN(dbg_0_dbg_uart_0_n_8_23));
	OAI211_X1_LVT dbg_0dbg_uart_0i_8_25 (.A(dbg_0_dbg_uart_0_n_8_11),.B(dbg_0_dbg_uart_0_n_8_14),.C1(dbg_0_dbg_uart_0_n_8_23),.C2(dbg_0_dbg_uart_0_n_8_24),.ZN(dbg_0_dbg_uart_0_uart_state_nxt_reg[0]));
	DFFR_X1_LVT dbg_0dbg_uart_0uart_state_reg___05F05b0___05F05d (.D(dbg_0_dbg_uart_0_uart_state_nxt_reg[0]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_23),.Q(dbg_0_dbg_uart_0_uart_state[0]),.QN());
	NOR3_X1_LVT dbg_0dbg_uart_0i_13_7 (.A1(dbg_0_dbg_uart_0_uart_state[0]),.A2(dbg_0_dbg_uart_0_uart_state[1]),.A3(dbg_0_dbg_uart_0_uart_state[2]),.ZN(dbg_0_dbg_uart_0_n_29));
	AND2_X1_LVT dbg_0dbg_uart_0i_17_0 (.A1(dbg_0_dbg_uart_0_n_29),.A2(dbg_0_dbg_uart_0_rxd_fe),.ZN(dbg_0_dbg_uart_0_n_33));
	OR2_X1_LVT dbg_0dbg_uart_0i_18_0 (.A1(dbg_0_dbg_uart_0_n_31),.A2(dbg_0_dbg_uart_0_n_33),.ZN(dbg_0_dbg_uart_0_n_34));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_busy_reg (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_34),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_32));
	DFFR_X1_LVT dbg_0dbg_uart_0sync_busy_reg (.D(dbg_0_dbg_uart_0_n_33),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_32),.Q(dbg_0_dbg_uart_0_sync_busy),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_22_0 (.A(dbg_0_dbg_uart_0_sync_busy),.ZN(dbg_0_dbg_uart_0_n_22_0));
	NAND2_X1_LVT dbg_0dbg_uart_0i_22_2 (.A1(dbg_0_dbg_uart_0_n_22_1),.A2(dbg_0_dbg_uart_0_n_22_0),.ZN(dbg_0_dbg_uart_0_n_76));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F14 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_50));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b3___05F05d (.D(dbg_0_dbg_uart_0_n_60),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_50),.Q(dbg_0_dbg_uart_0_bit_cnt_max[0]),.QN());
	HA_X1_LVT dbg_0dbg_uart_0i_21_3 (.A(dbg_0_dbg_uart_0_bit_cnt_max[0]),.B(dbg_0_dbg_uart_0_n_21_1),.CO(dbg_0_dbg_uart_0_n_21_2),.S(dbg_0_dbg_uart_0_n_60));
	HA_X1_LVT dbg_0dbg_uart_0i_21_4 (.A(dbg_0_dbg_uart_0_bit_cnt_max[1]),.B(dbg_0_dbg_uart_0_n_21_2),.CO(dbg_0_dbg_uart_0_n_21_3),.S(dbg_0_dbg_uart_0_n_61));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F13 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_49));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b4___05F05d (.D(dbg_0_dbg_uart_0_n_61),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_49),.Q(dbg_0_dbg_uart_0_bit_cnt_max[1]),.QN());
	XOR2_X1_LVT dbg_0dbg_uart_0i_29_0 (.A(dbg_0_dbg_uart_0_rxd_maj),.B(dbg_0_dbg_uart_0_rxd_maj_nxt),.Z(dbg_0_dbg_uart_0_n_29_0));
	AND2_X1_LVT dbg_0dbg_uart_0i_29_1 (.A1(dbg_0_dbg_uart_0_n_29_0),.A2(dbg_0_dbg_uart_0_rx_active),.ZN(dbg_0_dbg_uart_0_n_95));
	OR2_X1_LVT dbg_0dbg_uart_0i_28_0 (.A1(dbg_0_dbg_uart_0_txd_start),.A2(dbg_0_dbg_uart_0_xfer_bit_inc),.ZN(dbg_0_dbg_uart_0_n_94));
	INV_X1_LVT dbg_0dbg_uart_0i_30_1 (.A(dbg_0_dbg_uart_0_n_94),.ZN(dbg_0_dbg_uart_0_n_30_0));
	NOR2_X1_LVT dbg_0dbg_uart_0i_30_2 (.A1(dbg_0_dbg_uart_0_n_30_0),.A2(dbg_0_dbg_uart_0_n_95),.ZN(dbg_0_dbg_uart_0_n_97));
	INV_X1_LVT dbg_0dbg_uart_0i_27_0 (.A(dbg_0_dbg_uart_0_xfer_cnt[0]),.ZN(dbg_0_dbg_uart_0_n_78));
	NOR2_X1_LVT dbg_0dbg_uart_0i_30_0 (.A1(dbg_0_dbg_uart_0_n_94),.A2(dbg_0_dbg_uart_0_n_95),.ZN(dbg_0_dbg_uart_0_n_96));
	AOI222_X1_LVT dbg_0dbg_uart_0i_31_0 (.A1(dbg_0_dbg_uart_0_bit_cnt_max[1]),.A2(dbg_0_dbg_uart_0_n_95),.B1(dbg_0_dbg_uart_0_bit_cnt_max[0]),.B2(dbg_0_dbg_uart_0_n_97),.C1(dbg_0_dbg_uart_0_n_78),.C2(dbg_0_dbg_uart_0_n_96),.ZN(dbg_0_dbg_uart_0_n_31_0));
	INV_X1_LVT dbg_0dbg_uart_0i_31_1 (.A(dbg_0_dbg_uart_0_n_31_0),.ZN(dbg_0_dbg_uart_0_n_98));
	INV_X1_LVT dbg_0dbg_uart_0i_33_0 (.A(dbg_0_dbg_uart_0_n_94),.ZN(dbg_0_dbg_uart_0_n_33_0));
	INV_X1_LVT dbg_0dbg_uart_0i_33_1 (.A(dbg_0_dbg_uart_0_n_95),.ZN(dbg_0_dbg_uart_0_n_33_1));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_1 (.A(dbg_0_dbg_uart_0_xfer_cnt[1]),.B(dbg_0_dbg_uart_0_xfer_cnt[0]),.ZN(dbg_0_dbg_uart_0_n_79));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_2 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_79),.ZN(dbg_0_dbg_uart_0_n_31_1));
	INV_X1_LVT dbg_0dbg_uart_0i_31_3 (.A(dbg_0_dbg_uart_0_n_95),.ZN(dbg_0_dbg_uart_0_n_31_2));
	HA_X1_LVT dbg_0dbg_uart_0i_21_5 (.A(dbg_0_dbg_uart_0_bit_cnt_max[2]),.B(dbg_0_dbg_uart_0_n_21_3),.CO(dbg_0_dbg_uart_0_n_21_4),.S(dbg_0_dbg_uart_0_n_62));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F12 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_48));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b5___05F05d (.D(dbg_0_dbg_uart_0_n_62),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_48),.Q(dbg_0_dbg_uart_0_bit_cnt_max[2]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_4 (.A(dbg_0_dbg_uart_0_bit_cnt_max[2]),.ZN(dbg_0_dbg_uart_0_n_31_3));
	INV_X1_LVT dbg_0dbg_uart_0i_31_5 (.A(dbg_0_dbg_uart_0_bit_cnt_max[1]),.ZN(dbg_0_dbg_uart_0_n_31_4));
	INV_X1_LVT dbg_0dbg_uart_0i_31_6 (.A(dbg_0_dbg_uart_0_n_97),.ZN(dbg_0_dbg_uart_0_n_31_5));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_7 (.A(dbg_0_dbg_uart_0_n_31_1),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_3),.C1(dbg_0_dbg_uart_0_n_31_4),.C2(dbg_0_dbg_uart_0_n_31_5),.ZN(dbg_0_dbg_uart_0_n_99));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b1___05F05d (.D(dbg_0_dbg_uart_0_n_99),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[1]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_2 (.A1(dbg_0_dbg_uart_0_xfer_cnt[1]),.A2(dbg_0_dbg_uart_0_xfer_cnt[0]),.ZN(dbg_0_dbg_uart_0_n_27_0));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_3 (.A(dbg_0_dbg_uart_0_xfer_cnt[2]),.B(dbg_0_dbg_uart_0_n_27_0),.ZN(dbg_0_dbg_uart_0_n_80));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_8 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_80),.ZN(dbg_0_dbg_uart_0_n_31_6));
	HA_X1_LVT dbg_0dbg_uart_0i_21_6 (.A(dbg_0_dbg_uart_0_bit_cnt_max[3]),.B(dbg_0_dbg_uart_0_n_21_4),.CO(dbg_0_dbg_uart_0_n_21_5),.S(dbg_0_dbg_uart_0_n_63));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F11 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_47));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b6___05F05d (.D(dbg_0_dbg_uart_0_n_63),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_47),.Q(dbg_0_dbg_uart_0_bit_cnt_max[3]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_9 (.A(dbg_0_dbg_uart_0_bit_cnt_max[3]),.ZN(dbg_0_dbg_uart_0_n_31_7));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_10 (.A(dbg_0_dbg_uart_0_n_31_6),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_7),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_3),.ZN(dbg_0_dbg_uart_0_n_100));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b2___05F05d (.D(dbg_0_dbg_uart_0_n_100),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[2]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_4 (.A1(dbg_0_dbg_uart_0_xfer_cnt[2]),.A2(dbg_0_dbg_uart_0_n_27_0),.ZN(dbg_0_dbg_uart_0_n_27_1));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_5 (.A(dbg_0_dbg_uart_0_xfer_cnt[3]),.B(dbg_0_dbg_uart_0_n_27_1),.ZN(dbg_0_dbg_uart_0_n_81));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_11 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_81),.ZN(dbg_0_dbg_uart_0_n_31_8));
	HA_X1_LVT dbg_0dbg_uart_0i_21_7 (.A(dbg_0_dbg_uart_0_bit_cnt_max[4]),.B(dbg_0_dbg_uart_0_n_21_5),.CO(dbg_0_dbg_uart_0_n_21_6),.S(dbg_0_dbg_uart_0_n_64));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F10 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_46));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b7___05F05d (.D(dbg_0_dbg_uart_0_n_64),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_46),.Q(dbg_0_dbg_uart_0_bit_cnt_max[4]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_12 (.A(dbg_0_dbg_uart_0_bit_cnt_max[4]),.ZN(dbg_0_dbg_uart_0_n_31_9));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_13 (.A(dbg_0_dbg_uart_0_n_31_8),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_9),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_7),.ZN(dbg_0_dbg_uart_0_n_101));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b3___05F05d (.D(dbg_0_dbg_uart_0_n_101),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[3]),.QN());
	NOR4_X1_LVT dbg_0dbg_uart_0i_32_0 (.A1(dbg_0_dbg_uart_0_xfer_cnt[0]),.A2(dbg_0_dbg_uart_0_xfer_cnt[1]),.A3(dbg_0_dbg_uart_0_xfer_cnt[2]),.A4(dbg_0_dbg_uart_0_xfer_cnt[3]),.ZN(dbg_0_dbg_uart_0_n_32_0));
	OR2_X1_LVT dbg_0dbg_uart_0i_27_6 (.A1(dbg_0_dbg_uart_0_xfer_cnt[3]),.A2(dbg_0_dbg_uart_0_n_27_1),.ZN(dbg_0_dbg_uart_0_n_27_2));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_7 (.A(dbg_0_dbg_uart_0_xfer_cnt[4]),.B(dbg_0_dbg_uart_0_n_27_2),.ZN(dbg_0_dbg_uart_0_n_82));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_14 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_82),.ZN(dbg_0_dbg_uart_0_n_31_10));
	HA_X1_LVT dbg_0dbg_uart_0i_21_8 (.A(dbg_0_dbg_uart_0_bit_cnt_max[5]),.B(dbg_0_dbg_uart_0_n_21_6),.CO(dbg_0_dbg_uart_0_n_21_7),.S(dbg_0_dbg_uart_0_n_65));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F9 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_45));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b8___05F05d (.D(dbg_0_dbg_uart_0_n_65),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_45),.Q(dbg_0_dbg_uart_0_bit_cnt_max[5]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_15 (.A(dbg_0_dbg_uart_0_bit_cnt_max[5]),.ZN(dbg_0_dbg_uart_0_n_31_11));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_16 (.A(dbg_0_dbg_uart_0_n_31_10),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_11),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_9),.ZN(dbg_0_dbg_uart_0_n_102));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b4___05F05d (.D(dbg_0_dbg_uart_0_n_102),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[4]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_8 (.A1(dbg_0_dbg_uart_0_xfer_cnt[4]),.A2(dbg_0_dbg_uart_0_n_27_2),.ZN(dbg_0_dbg_uart_0_n_27_3));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_9 (.A(dbg_0_dbg_uart_0_xfer_cnt[5]),.B(dbg_0_dbg_uart_0_n_27_3),.ZN(dbg_0_dbg_uart_0_n_83));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_17 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_83),.ZN(dbg_0_dbg_uart_0_n_31_12));
	HA_X1_LVT dbg_0dbg_uart_0i_21_9 (.A(dbg_0_dbg_uart_0_bit_cnt_max[6]),.B(dbg_0_dbg_uart_0_n_21_7),.CO(dbg_0_dbg_uart_0_n_21_8),.S(dbg_0_dbg_uart_0_n_66));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F8 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_44));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b9___05F05d (.D(dbg_0_dbg_uart_0_n_66),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_44),.Q(dbg_0_dbg_uart_0_bit_cnt_max[6]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_18 (.A(dbg_0_dbg_uart_0_bit_cnt_max[6]),.ZN(dbg_0_dbg_uart_0_n_31_13));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_19 (.A(dbg_0_dbg_uart_0_n_31_12),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_13),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_11),.ZN(dbg_0_dbg_uart_0_n_103));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b5___05F05d (.D(dbg_0_dbg_uart_0_n_103),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[5]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_10 (.A1(dbg_0_dbg_uart_0_xfer_cnt[5]),.A2(dbg_0_dbg_uart_0_n_27_3),.ZN(dbg_0_dbg_uart_0_n_27_4));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_11 (.A(dbg_0_dbg_uart_0_xfer_cnt[6]),.B(dbg_0_dbg_uart_0_n_27_4),.ZN(dbg_0_dbg_uart_0_n_84));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_20 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_84),.ZN(dbg_0_dbg_uart_0_n_31_14));
	HA_X1_LVT dbg_0dbg_uart_0i_21_10 (.A(dbg_0_dbg_uart_0_bit_cnt_max[7]),.B(dbg_0_dbg_uart_0_n_21_8),.CO(dbg_0_dbg_uart_0_n_21_9),.S(dbg_0_dbg_uart_0_n_67));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F7 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_43));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b10___05F05d (.D(dbg_0_dbg_uart_0_n_67),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_43),.Q(dbg_0_dbg_uart_0_bit_cnt_max[7]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_21 (.A(dbg_0_dbg_uart_0_bit_cnt_max[7]),.ZN(dbg_0_dbg_uart_0_n_31_15));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_22 (.A(dbg_0_dbg_uart_0_n_31_14),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_15),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_13),.ZN(dbg_0_dbg_uart_0_n_104));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b6___05F05d (.D(dbg_0_dbg_uart_0_n_104),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[6]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_12 (.A1(dbg_0_dbg_uart_0_xfer_cnt[6]),.A2(dbg_0_dbg_uart_0_n_27_4),.ZN(dbg_0_dbg_uart_0_n_27_5));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_13 (.A(dbg_0_dbg_uart_0_xfer_cnt[7]),.B(dbg_0_dbg_uart_0_n_27_5),.ZN(dbg_0_dbg_uart_0_n_85));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_23 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_85),.ZN(dbg_0_dbg_uart_0_n_31_16));
	HA_X1_LVT dbg_0dbg_uart_0i_21_11 (.A(dbg_0_dbg_uart_0_bit_cnt_max[8]),.B(dbg_0_dbg_uart_0_n_21_9),.CO(dbg_0_dbg_uart_0_n_21_10),.S(dbg_0_dbg_uart_0_n_68));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F6 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_42));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b11___05F05d (.D(dbg_0_dbg_uart_0_n_68),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_42),.Q(dbg_0_dbg_uart_0_bit_cnt_max[8]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_24 (.A(dbg_0_dbg_uart_0_bit_cnt_max[8]),.ZN(dbg_0_dbg_uart_0_n_31_17));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_25 (.A(dbg_0_dbg_uart_0_n_31_16),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_17),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_15),.ZN(dbg_0_dbg_uart_0_n_105));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b7___05F05d (.D(dbg_0_dbg_uart_0_n_105),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[7]),.QN());
	NOR4_X1_LVT dbg_0dbg_uart_0i_32_1 (.A1(dbg_0_dbg_uart_0_xfer_cnt[4]),.A2(dbg_0_dbg_uart_0_xfer_cnt[5]),.A3(dbg_0_dbg_uart_0_xfer_cnt[6]),.A4(dbg_0_dbg_uart_0_xfer_cnt[7]),.ZN(dbg_0_dbg_uart_0_n_32_1));
	OR2_X1_LVT dbg_0dbg_uart_0i_27_14 (.A1(dbg_0_dbg_uart_0_xfer_cnt[7]),.A2(dbg_0_dbg_uart_0_n_27_5),.ZN(dbg_0_dbg_uart_0_n_27_6));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_15 (.A(dbg_0_dbg_uart_0_xfer_cnt[8]),.B(dbg_0_dbg_uart_0_n_27_6),.ZN(dbg_0_dbg_uart_0_n_86));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_26 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_86),.ZN(dbg_0_dbg_uart_0_n_31_18));
	HA_X1_LVT dbg_0dbg_uart_0i_21_12 (.A(dbg_0_dbg_uart_0_bit_cnt_max[9]),.B(dbg_0_dbg_uart_0_n_21_10),.CO(dbg_0_dbg_uart_0_n_21_11),.S(dbg_0_dbg_uart_0_n_69));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F5 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_41));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b12___05F05d (.D(dbg_0_dbg_uart_0_n_69),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_41),.Q(dbg_0_dbg_uart_0_bit_cnt_max[9]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_27 (.A(dbg_0_dbg_uart_0_bit_cnt_max[9]),.ZN(dbg_0_dbg_uart_0_n_31_19));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_28 (.A(dbg_0_dbg_uart_0_n_31_18),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_19),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_17),.ZN(dbg_0_dbg_uart_0_n_106));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b8___05F05d (.D(dbg_0_dbg_uart_0_n_106),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[8]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_16 (.A1(dbg_0_dbg_uart_0_xfer_cnt[8]),.A2(dbg_0_dbg_uart_0_n_27_6),.ZN(dbg_0_dbg_uart_0_n_27_7));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_17 (.A(dbg_0_dbg_uart_0_xfer_cnt[9]),.B(dbg_0_dbg_uart_0_n_27_7),.ZN(dbg_0_dbg_uart_0_n_87));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_29 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_87),.ZN(dbg_0_dbg_uart_0_n_31_20));
	HA_X1_LVT dbg_0dbg_uart_0i_21_13 (.A(dbg_0_dbg_uart_0_bit_cnt_max[10]),.B(dbg_0_dbg_uart_0_n_21_11),.CO(dbg_0_dbg_uart_0_n_21_12),.S(dbg_0_dbg_uart_0_n_70));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F4 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_40));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b13___05F05d (.D(dbg_0_dbg_uart_0_n_70),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_40),.Q(dbg_0_dbg_uart_0_bit_cnt_max[10]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_30 (.A(dbg_0_dbg_uart_0_bit_cnt_max[10]),.ZN(dbg_0_dbg_uart_0_n_31_21));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_31 (.A(dbg_0_dbg_uart_0_n_31_20),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_21),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_19),.ZN(dbg_0_dbg_uart_0_n_107));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b9___05F05d (.D(dbg_0_dbg_uart_0_n_107),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[9]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_18 (.A1(dbg_0_dbg_uart_0_xfer_cnt[9]),.A2(dbg_0_dbg_uart_0_n_27_7),.ZN(dbg_0_dbg_uart_0_n_27_8));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_19 (.A(dbg_0_dbg_uart_0_xfer_cnt[10]),.B(dbg_0_dbg_uart_0_n_27_8),.ZN(dbg_0_dbg_uart_0_n_88));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_32 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_88),.ZN(dbg_0_dbg_uart_0_n_31_22));
	HA_X1_LVT dbg_0dbg_uart_0i_21_14 (.A(dbg_0_dbg_uart_0_bit_cnt_max[11]),.B(dbg_0_dbg_uart_0_n_21_12),.CO(dbg_0_dbg_uart_0_n_21_13),.S(dbg_0_dbg_uart_0_n_71));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F3 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_39));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b14___05F05d (.D(dbg_0_dbg_uart_0_n_71),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_39),.Q(dbg_0_dbg_uart_0_bit_cnt_max[11]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_33 (.A(dbg_0_dbg_uart_0_bit_cnt_max[11]),.ZN(dbg_0_dbg_uart_0_n_31_23));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_34 (.A(dbg_0_dbg_uart_0_n_31_22),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_23),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_21),.ZN(dbg_0_dbg_uart_0_n_108));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b10___05F05d (.D(dbg_0_dbg_uart_0_n_108),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[10]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_20 (.A1(dbg_0_dbg_uart_0_xfer_cnt[10]),.A2(dbg_0_dbg_uart_0_n_27_8),.ZN(dbg_0_dbg_uart_0_n_27_9));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_21 (.A(dbg_0_dbg_uart_0_xfer_cnt[11]),.B(dbg_0_dbg_uart_0_n_27_9),.ZN(dbg_0_dbg_uart_0_n_89));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_35 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_89),.ZN(dbg_0_dbg_uart_0_n_31_24));
	HA_X1_LVT dbg_0dbg_uart_0i_21_15 (.A(dbg_0_dbg_uart_0_bit_cnt_max[12]),.B(dbg_0_dbg_uart_0_n_21_13),.CO(dbg_0_dbg_uart_0_n_21_14),.S(dbg_0_dbg_uart_0_n_72));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F2 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_38));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b15___05F05d (.D(dbg_0_dbg_uart_0_n_72),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_38),.Q(dbg_0_dbg_uart_0_bit_cnt_max[12]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_36 (.A(dbg_0_dbg_uart_0_bit_cnt_max[12]),.ZN(dbg_0_dbg_uart_0_n_31_25));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_37 (.A(dbg_0_dbg_uart_0_n_31_24),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_25),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_23),.ZN(dbg_0_dbg_uart_0_n_109));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b11___05F05d (.D(dbg_0_dbg_uart_0_n_109),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[11]),.QN());
	NOR4_X1_LVT dbg_0dbg_uart_0i_32_2 (.A1(dbg_0_dbg_uart_0_xfer_cnt[8]),.A2(dbg_0_dbg_uart_0_xfer_cnt[9]),.A3(dbg_0_dbg_uart_0_xfer_cnt[10]),.A4(dbg_0_dbg_uart_0_xfer_cnt[11]),.ZN(dbg_0_dbg_uart_0_n_32_2));
	OR2_X1_LVT dbg_0dbg_uart_0i_27_22 (.A1(dbg_0_dbg_uart_0_xfer_cnt[11]),.A2(dbg_0_dbg_uart_0_n_27_9),.ZN(dbg_0_dbg_uart_0_n_27_10));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_23 (.A(dbg_0_dbg_uart_0_xfer_cnt[12]),.B(dbg_0_dbg_uart_0_n_27_10),.ZN(dbg_0_dbg_uart_0_n_90));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_38 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_90),.ZN(dbg_0_dbg_uart_0_n_31_26));
	HA_X1_LVT dbg_0dbg_uart_0i_21_16 (.A(dbg_0_dbg_uart_0_bit_cnt_max[13]),.B(dbg_0_dbg_uart_0_n_21_14),.CO(dbg_0_dbg_uart_0_n_21_15),.S(dbg_0_dbg_uart_0_n_73));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F1 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_37));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b16___05F05d (.D(dbg_0_dbg_uart_0_n_73),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_37),.Q(dbg_0_dbg_uart_0_bit_cnt_max[13]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_39 (.A(dbg_0_dbg_uart_0_bit_cnt_max[13]),.ZN(dbg_0_dbg_uart_0_n_31_27));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_40 (.A(dbg_0_dbg_uart_0_n_31_26),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_27),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_25),.ZN(dbg_0_dbg_uart_0_n_110));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b12___05F05d (.D(dbg_0_dbg_uart_0_n_110),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[12]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_24 (.A1(dbg_0_dbg_uart_0_xfer_cnt[12]),.A2(dbg_0_dbg_uart_0_n_27_10),.ZN(dbg_0_dbg_uart_0_n_27_11));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_25 (.A(dbg_0_dbg_uart_0_xfer_cnt[13]),.B(dbg_0_dbg_uart_0_n_27_11),.ZN(dbg_0_dbg_uart_0_n_91));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_41 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_91),.ZN(dbg_0_dbg_uart_0_n_31_28));
	HA_X1_LVT dbg_0dbg_uart_0i_21_17 (.A(dbg_0_dbg_uart_0_bit_cnt_max[14]),.B(dbg_0_dbg_uart_0_n_21_15),.CO(dbg_0_dbg_uart_0_n_21_16),.S(dbg_0_dbg_uart_0_n_74));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg___05F_05F0 (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_36));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b17___05F05d (.D(dbg_0_dbg_uart_0_n_74),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_36),.Q(dbg_0_dbg_uart_0_bit_cnt_max[14]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_42 (.A(dbg_0_dbg_uart_0_bit_cnt_max[14]),.ZN(dbg_0_dbg_uart_0_n_31_29));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_43 (.A(dbg_0_dbg_uart_0_n_31_28),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_29),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_27),.ZN(dbg_0_dbg_uart_0_n_111));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b13___05F05d (.D(dbg_0_dbg_uart_0_n_111),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[13]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_26 (.A1(dbg_0_dbg_uart_0_xfer_cnt[13]),.A2(dbg_0_dbg_uart_0_n_27_11),.ZN(dbg_0_dbg_uart_0_n_27_12));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_27 (.A(dbg_0_dbg_uart_0_xfer_cnt[14]),.B(dbg_0_dbg_uart_0_n_27_12),.ZN(dbg_0_dbg_uart_0_n_92));
	NAND2_X1_LVT dbg_0dbg_uart_0i_31_44 (.A1(dbg_0_dbg_uart_0_n_96),.A2(dbg_0_dbg_uart_0_n_92),.ZN(dbg_0_dbg_uart_0_n_31_30));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_21_18 (.A(dbg_0_dbg_uart_0_bit_cnt_max[15]),.B(dbg_0_dbg_uart_0_n_21_16),.ZN(dbg_0_dbg_uart_0_n_21_17));
	INV_X1_LVT dbg_0dbg_uart_0i_21_19 (.A(dbg_0_dbg_uart_0_n_21_17),.ZN(dbg_0_dbg_uart_0_n_75));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_sync_cnt_reg (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_76),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_35));
	DFFS_X1_LVT dbg_0dbg_uart_0sync_cnt_reg___05F05b18___05F05d (.D(dbg_0_dbg_uart_0_n_75),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_35),.Q(dbg_0_dbg_uart_0_bit_cnt_max[15]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_31_45 (.A(dbg_0_dbg_uart_0_bit_cnt_max[15]),.ZN(dbg_0_dbg_uart_0_n_31_31));
	OAI221_X1_LVT dbg_0dbg_uart_0i_31_46 (.A(dbg_0_dbg_uart_0_n_31_30),.B1(dbg_0_dbg_uart_0_n_31_2),.B2(dbg_0_dbg_uart_0_n_31_31),.C1(dbg_0_dbg_uart_0_n_31_5),.C2(dbg_0_dbg_uart_0_n_31_29),.ZN(dbg_0_dbg_uart_0_n_112));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b14___05F05d (.D(dbg_0_dbg_uart_0_n_112),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[14]),.QN());
	OR2_X1_LVT dbg_0dbg_uart_0i_27_28 (.A1(dbg_0_dbg_uart_0_xfer_cnt[14]),.A2(dbg_0_dbg_uart_0_n_27_12),.ZN(dbg_0_dbg_uart_0_n_27_13));
	XNOR2_X1_LVT dbg_0dbg_uart_0i_27_29 (.A(dbg_0_dbg_uart_0_xfer_cnt[15]),.B(dbg_0_dbg_uart_0_n_27_13),.ZN(dbg_0_dbg_uart_0_n_93));
	AOI22_X1_LVT dbg_0dbg_uart_0i_31_47 (.A1(dbg_0_dbg_uart_0_n_97),.A2(dbg_0_dbg_uart_0_bit_cnt_max[15]),.B1(dbg_0_dbg_uart_0_n_96),.B2(dbg_0_dbg_uart_0_n_93),.ZN(dbg_0_dbg_uart_0_n_31_32));
	INV_X1_LVT dbg_0dbg_uart_0i_31_48 (.A(dbg_0_dbg_uart_0_n_31_32),.ZN(dbg_0_dbg_uart_0_n_113));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b15___05F05d (.D(dbg_0_dbg_uart_0_n_113),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[15]),.QN());
	NOR4_X1_LVT dbg_0dbg_uart_0i_32_3 (.A1(dbg_0_dbg_uart_0_xfer_cnt[12]),.A2(dbg_0_dbg_uart_0_xfer_cnt[13]),.A3(dbg_0_dbg_uart_0_xfer_cnt[14]),.A4(dbg_0_dbg_uart_0_xfer_cnt[15]),.ZN(dbg_0_dbg_uart_0_n_32_3));
	NAND4_X1_LVT dbg_0dbg_uart_0i_32_4 (.A1(dbg_0_dbg_uart_0_n_32_0),.A2(dbg_0_dbg_uart_0_n_32_1),.A3(dbg_0_dbg_uart_0_n_32_2),.A4(dbg_0_dbg_uart_0_n_32_3),.ZN(dbg_0_dbg_uart_0_n_114));
	NAND3_X1_LVT dbg_0dbg_uart_0i_33_2 (.A1(dbg_0_dbg_uart_0_n_33_0),.A2(dbg_0_dbg_uart_0_n_33_1),.A3(dbg_0_dbg_uart_0_n_114),.ZN(dbg_0_dbg_uart_0_n_33_2));
	NAND3_X1_LVT dbg_0dbg_uart_0i_33_3 (.A1(dbg_0_dbg_uart_0_n_33_2),.A2(dbg_0_dbg_uart_0_n_33_0),.A3(dbg_0_dbg_uart_0_n_33_1),.ZN(dbg_0_dbg_uart_0_n_115));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_xfer_cnt_reg (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_115),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_77));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_cnt_reg___05F05b0___05F05d (.D(dbg_0_dbg_uart_0_n_98),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_77),.Q(dbg_0_dbg_uart_0_xfer_cnt[0]),.QN());
	NOR4_X1_LVT dbg_0dbg_uart_0i_35_0 (.A1(dbg_0_dbg_uart_0_xfer_cnt[0]),.A2(dbg_0_dbg_uart_0_xfer_cnt[1]),.A3(dbg_0_dbg_uart_0_xfer_cnt[2]),.A4(dbg_0_dbg_uart_0_xfer_cnt[3]),.ZN(dbg_0_dbg_uart_0_n_35_0));
	NOR4_X1_LVT dbg_0dbg_uart_0i_35_1 (.A1(dbg_0_dbg_uart_0_xfer_cnt[4]),.A2(dbg_0_dbg_uart_0_xfer_cnt[5]),.A3(dbg_0_dbg_uart_0_xfer_cnt[6]),.A4(dbg_0_dbg_uart_0_xfer_cnt[7]),.ZN(dbg_0_dbg_uart_0_n_35_1));
	NOR4_X1_LVT dbg_0dbg_uart_0i_35_2 (.A1(dbg_0_dbg_uart_0_xfer_cnt[8]),.A2(dbg_0_dbg_uart_0_xfer_cnt[9]),.A3(dbg_0_dbg_uart_0_xfer_cnt[10]),.A4(dbg_0_dbg_uart_0_xfer_cnt[11]),.ZN(dbg_0_dbg_uart_0_n_35_2));
	NOR4_X1_LVT dbg_0dbg_uart_0i_35_3 (.A1(dbg_0_dbg_uart_0_xfer_cnt[12]),.A2(dbg_0_dbg_uart_0_xfer_cnt[13]),.A3(dbg_0_dbg_uart_0_xfer_cnt[14]),.A4(dbg_0_dbg_uart_0_xfer_cnt[15]),.ZN(dbg_0_dbg_uart_0_n_35_3));
	NAND4_X1_LVT dbg_0dbg_uart_0i_35_4 (.A1(dbg_0_dbg_uart_0_n_35_0),.A2(dbg_0_dbg_uart_0_n_35_1),.A3(dbg_0_dbg_uart_0_n_35_2),.A4(dbg_0_dbg_uart_0_n_35_3),.ZN(dbg_0_dbg_uart_0_n_35_4));
	NOR4_X1_LVT dbg_0dbg_uart_0i_35_5 (.A1(dbg_0_dbg_uart_0_xfer_bit[0]),.A2(dbg_0_dbg_uart_0_xfer_bit[1]),.A3(dbg_0_dbg_uart_0_xfer_bit[2]),.A4(dbg_0_dbg_uart_0_xfer_bit[3]),.ZN(dbg_0_dbg_uart_0_n_35_5));
	NOR2_X1_LVT dbg_0dbg_uart_0i_35_6 (.A1(dbg_0_dbg_uart_0_n_35_4),.A2(dbg_0_dbg_uart_0_n_35_5),.ZN(dbg_0_dbg_uart_0_xfer_bit_inc));
	INV_X1_LVT dbg_0dbg_uart_0i_5_1 (.A(dbg_0_dbg_uart_0_xfer_bit_inc),.ZN(dbg_0_dbg_uart_0_n_5_1));
	INV_X1_LVT dbg_0dbg_uart_0i_5_0 (.A(dbg_0_dbg_rd_rdy),.ZN(dbg_0_dbg_uart_0_n_5_0));
	NAND2_X1_LVT dbg_0dbg_uart_0i_5_2 (.A1(dbg_0_dbg_uart_0_n_5_1),.A2(dbg_0_dbg_uart_0_n_5_0),.ZN(dbg_0_dbg_uart_0_n_21));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_xfer_buf_reg (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_21),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_0));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b19___05F05d (.D(dbg_0_dbg_uart_0_n_19),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[0]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_34 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[15]),.ZN(dbg_0_dbg_uart_0_n_4_17));
	INV_X1_LVT dbg_0dbg_uart_0i_4_35 (.A(dbg_0_dbg_uart_0_n_4_17),.ZN(dbg_0_dbg_uart_0_n_18));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b18___05F05d (.D(dbg_0_dbg_uart_0_n_18),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[0]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_32 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[14]),.ZN(dbg_0_dbg_uart_0_n_4_16));
	INV_X1_LVT dbg_0dbg_uart_0i_4_33 (.A(dbg_0_dbg_uart_0_n_4_16),.ZN(dbg_0_dbg_uart_0_n_17));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b17___05F05d (.D(dbg_0_dbg_uart_0_n_17),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[0]),.QN());
	AND2_X1_LVT dbg_0dbg_uart_0i_45_0 (.A1(dbg_0_dbg_uart_0_n_27),.A2(dbg_0_dbg_uart_0_xfer_done),.ZN(dbg_0_dbg_uart_0_cmd_valid));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_dbg_addr_reg (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_cmd_valid),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_129));
	DFFR_X1_LVT dbg_0dbg_uart_0dbg_addr_reg___05F05b5___05F05d (.D(dbg_0_dbg_uart_0_xfer_buf[0]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_129),.Q(dbg_0_dbg_addr[5]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_30 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[13]),.ZN(dbg_0_dbg_uart_0_n_4_15));
	INV_X1_LVT dbg_0dbg_uart_0i_4_31 (.A(dbg_0_dbg_uart_0_n_4_15),.ZN(dbg_0_dbg_uart_0_n_16));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b16___05F05d (.D(dbg_0_dbg_uart_0_n_16),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[0]),.QN());
	DFFR_X1_LVT dbg_0dbg_uart_0dbg_addr_reg___05F05b4___05F05d (.D(dbg_0_dbg_uart_0_xfer_buf[0]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_129),.Q(dbg_0_dbg_addr[4]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_28 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[12]),.ZN(dbg_0_dbg_uart_0_n_4_14));
	INV_X1_LVT dbg_0dbg_uart_0i_4_29 (.A(dbg_0_dbg_uart_0_n_4_14),.ZN(dbg_0_dbg_uart_0_n_15));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b15___05F05d (.D(dbg_0_dbg_uart_0_n_15),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[15]),.QN());
	DFFR_X1_LVT dbg_0dbg_uart_0dbg_addr_reg___05F05b3___05F05d (.D(dbg_0_dbg_uart_0_xfer_buf[15]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_129),.Q(dbg_0_dbg_addr[3]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_26 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[15]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[11]),.ZN(dbg_0_dbg_uart_0_n_4_13));
	INV_X1_LVT dbg_0dbg_uart_0i_4_27 (.A(dbg_0_dbg_uart_0_n_4_13),.ZN(dbg_0_dbg_uart_0_n_14));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b14___05F05d (.D(dbg_0_dbg_uart_0_n_14),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[14]),.QN());
	DFFR_X1_LVT dbg_0dbg_uart_0dbg_addr_reg___05F05b2___05F05d (.D(dbg_0_dbg_uart_0_xfer_buf[14]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_129),.Q(dbg_0_dbg_addr[2]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_24 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[14]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[10]),.ZN(dbg_0_dbg_uart_0_n_4_12));
	INV_X1_LVT dbg_0dbg_uart_0i_4_25 (.A(dbg_0_dbg_uart_0_n_4_12),.ZN(dbg_0_dbg_uart_0_n_13));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b13___05F05d (.D(dbg_0_dbg_uart_0_n_13),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[13]),.QN());
	DFFR_X1_LVT dbg_0dbg_uart_0dbg_addr_reg___05F05b1___05F05d (.D(dbg_0_dbg_uart_0_xfer_buf[13]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_129),.Q(dbg_0_dbg_addr[1]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_22 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[13]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[9]),.ZN(dbg_0_dbg_uart_0_n_4_11));
	INV_X1_LVT dbg_0dbg_uart_0i_4_23 (.A(dbg_0_dbg_uart_0_n_4_11),.ZN(dbg_0_dbg_uart_0_n_12));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b12___05F05d (.D(dbg_0_dbg_uart_0_n_12),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[12]),.QN());
	DFFR_X1_LVT dbg_0dbg_uart_0dbg_addr_reg___05F05b0___05F05d (.D(dbg_0_dbg_uart_0_xfer_buf[12]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_129),.Q(dbg_0_dbg_addr[0]),.QN());
	INV_X1_LVT dbg_0dbg_uart_0i_49_0 (.A(dbg_0_mem_burst),.ZN(dbg_0_dbg_uart_0_n_49_0));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_dbg_bw_reg (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_cmd_valid),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_131));
	DFFR_X1_LVT dbg_0dbg_uart_0dbg_bw_reg (.D(dbg_0_dbg_uart_0_xfer_buf[0]),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_131),.Q(dbg_0_dbg_uart_0_dbg_bw),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_49_1 (.A1(dbg_0_dbg_uart_0_n_49_0),.A2(dbg_0_dbg_uart_0_dbg_bw),.B1(dbg_0_mem_ctl[2]),.B2(dbg_0_mem_burst),.ZN(dbg_0_dbg_uart_0_n_49_1));
	AND2_X1_LVT dbg_0dbg_uart_0i_49_26 (.A1(dbg_0_dbg_uart_0_n_49_1),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.ZN(dbg_0_dbg_din[15]));
	AND2_X1_LVT dbg_0dbg_uart_0i_49_25 (.A1(dbg_0_dbg_uart_0_n_49_1),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.ZN(dbg_0_dbg_din[14]));
	AND2_X1_LVT dbg_0dbg_uart_0i_49_24 (.A1(dbg_0_dbg_uart_0_n_49_1),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.ZN(dbg_0_dbg_din[13]));
	AND2_X1_LVT dbg_0dbg_uart_0i_49_23 (.A1(dbg_0_dbg_uart_0_n_49_1),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.ZN(dbg_0_dbg_din[12]));
	AND2_X1_LVT dbg_0dbg_uart_0i_49_22 (.A1(dbg_0_dbg_uart_0_n_49_1),.A2(dbg_0_dbg_uart_0_xfer_buf[15]),.ZN(dbg_0_dbg_din[11]));
	AND2_X1_LVT dbg_0dbg_uart_0i_49_21 (.A1(dbg_0_dbg_uart_0_n_49_1),.A2(dbg_0_dbg_uart_0_xfer_buf[14]),.ZN(dbg_0_dbg_din[10]));
	AND2_X1_LVT dbg_0dbg_uart_0i_49_20 (.A1(dbg_0_dbg_uart_0_n_49_1),.A2(dbg_0_dbg_uart_0_xfer_buf[13]),.ZN(dbg_0_dbg_din[9]));
	AND2_X1_LVT dbg_0dbg_uart_0i_49_19 (.A1(dbg_0_dbg_uart_0_n_49_1),.A2(dbg_0_dbg_uart_0_xfer_buf[12]),.ZN(dbg_0_dbg_din[8]));
	INV_X1_LVT dbg_0dbg_uart_0i_49_2 (.A(dbg_0_dbg_uart_0_n_49_1),.ZN(dbg_0_dbg_uart_0_n_49_2));
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_20 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[12]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[8]),.ZN(dbg_0_dbg_uart_0_n_4_10));
	INV_X1_LVT dbg_0dbg_uart_0i_4_21 (.A(dbg_0_dbg_uart_0_n_4_10),.ZN(dbg_0_dbg_uart_0_n_11));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b11___05F05d (.D(dbg_0_dbg_uart_0_n_11),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[11]),.QN());
	AND2_X1_LVT dbg_0dbg_uart_0i_4_19 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[11]),.ZN(dbg_0_dbg_uart_0_n_10));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b10___05F05d (.D(dbg_0_dbg_uart_0_n_10),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[10]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_49_17 (.A1(dbg_0_dbg_uart_0_n_49_2),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.B1(dbg_0_dbg_uart_0_n_49_1),.B2(dbg_0_dbg_uart_0_xfer_buf[10]),.ZN(dbg_0_dbg_uart_0_n_49_10));
	INV_X1_LVT dbg_0dbg_uart_0i_49_18 (.A(dbg_0_dbg_uart_0_n_49_10),.ZN(dbg_0_dbg_din[7]));
	INV_X1_LVT dbg_0dbg_uart_0i_4_18 (.A(dbg_0_dbg_uart_0_xfer_buf[10]),.ZN(dbg_0_dbg_uart_0_n_4_9));
	NAND2_X1_LVT dbg_0dbg_uart_0i_4_38 (.A1(dbg_0_dbg_uart_0_n_4_9),.A2(dbg_0_dbg_uart_0_n_4_0),.ZN(dbg_0_dbg_uart_0_n_20));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b9___05F05d (.D(dbg_0_dbg_uart_0_n_20),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[9]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_49_15 (.A1(dbg_0_dbg_uart_0_n_49_2),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.B1(dbg_0_dbg_uart_0_n_49_1),.B2(dbg_0_dbg_uart_0_xfer_buf[9]),.ZN(dbg_0_dbg_uart_0_n_49_9));
	INV_X1_LVT dbg_0dbg_uart_0i_49_16 (.A(dbg_0_dbg_uart_0_n_49_9),.ZN(dbg_0_dbg_din[6]));
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_16 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[9]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[7]),.ZN(dbg_0_dbg_uart_0_n_4_8));
	INV_X1_LVT dbg_0dbg_uart_0i_4_17 (.A(dbg_0_dbg_uart_0_n_4_8),.ZN(dbg_0_dbg_uart_0_n_9));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b8___05F05d (.D(dbg_0_dbg_uart_0_n_9),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[8]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_49_13 (.A1(dbg_0_dbg_uart_0_n_49_2),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.B1(dbg_0_dbg_uart_0_n_49_1),.B2(dbg_0_dbg_uart_0_xfer_buf[8]),.ZN(dbg_0_dbg_uart_0_n_49_8));
	INV_X1_LVT dbg_0dbg_uart_0i_49_14 (.A(dbg_0_dbg_uart_0_n_49_8),.ZN(dbg_0_dbg_din[5]));
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_14 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[8]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[6]),.ZN(dbg_0_dbg_uart_0_n_4_7));
	INV_X1_LVT dbg_0dbg_uart_0i_4_15 (.A(dbg_0_dbg_uart_0_n_4_7),.ZN(dbg_0_dbg_uart_0_n_8));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b7___05F05d (.D(dbg_0_dbg_uart_0_n_8),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[7]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_49_11 (.A1(dbg_0_dbg_uart_0_n_49_2),.A2(dbg_0_dbg_uart_0_xfer_buf[0]),.B1(dbg_0_dbg_uart_0_n_49_1),.B2(dbg_0_dbg_uart_0_xfer_buf[7]),.ZN(dbg_0_dbg_uart_0_n_49_7));
	INV_X1_LVT dbg_0dbg_uart_0i_49_12 (.A(dbg_0_dbg_uart_0_n_49_7),.ZN(dbg_0_dbg_din[4]));
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_12 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[7]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[5]),.ZN(dbg_0_dbg_uart_0_n_4_6));
	INV_X1_LVT dbg_0dbg_uart_0i_4_13 (.A(dbg_0_dbg_uart_0_n_4_6),.ZN(dbg_0_dbg_uart_0_n_7));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b6___05F05d (.D(dbg_0_dbg_uart_0_n_7),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[6]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_49_9 (.A1(dbg_0_dbg_uart_0_n_49_2),.A2(dbg_0_dbg_uart_0_xfer_buf[15]),.B1(dbg_0_dbg_uart_0_n_49_1),.B2(dbg_0_dbg_uart_0_xfer_buf[6]),.ZN(dbg_0_dbg_uart_0_n_49_6));
	INV_X1_LVT dbg_0dbg_uart_0i_49_10 (.A(dbg_0_dbg_uart_0_n_49_6),.ZN(dbg_0_dbg_din[3]));
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_10 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[6]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[4]),.ZN(dbg_0_dbg_uart_0_n_4_5));
	INV_X1_LVT dbg_0dbg_uart_0i_4_11 (.A(dbg_0_dbg_uart_0_n_4_5),.ZN(dbg_0_dbg_uart_0_n_6));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b5___05F05d (.D(dbg_0_dbg_uart_0_n_6),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[5]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_49_7 (.A1(dbg_0_dbg_uart_0_n_49_2),.A2(dbg_0_dbg_uart_0_xfer_buf[14]),.B1(dbg_0_dbg_uart_0_n_49_1),.B2(dbg_0_dbg_uart_0_xfer_buf[5]),.ZN(dbg_0_dbg_uart_0_n_49_5));
	INV_X1_LVT dbg_0dbg_uart_0i_49_8 (.A(dbg_0_dbg_uart_0_n_49_5),.ZN(dbg_0_dbg_din[2]));
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_8 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[5]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[3]),.ZN(dbg_0_dbg_uart_0_n_4_4));
	INV_X1_LVT dbg_0dbg_uart_0i_4_9 (.A(dbg_0_dbg_uart_0_n_4_4),.ZN(dbg_0_dbg_uart_0_n_5));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b4___05F05d (.D(dbg_0_dbg_uart_0_n_5),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[4]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_49_5 (.A1(dbg_0_dbg_uart_0_n_49_2),.A2(dbg_0_dbg_uart_0_xfer_buf[13]),.B1(dbg_0_dbg_uart_0_n_49_1),.B2(dbg_0_dbg_uart_0_xfer_buf[4]),.ZN(dbg_0_dbg_uart_0_n_49_4));
	INV_X1_LVT dbg_0dbg_uart_0i_49_6 (.A(dbg_0_dbg_uart_0_n_49_4),.ZN(dbg_0_dbg_din[1]));
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_6 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[4]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[2]),.ZN(dbg_0_dbg_uart_0_n_4_3));
	INV_X1_LVT dbg_0dbg_uart_0i_4_7 (.A(dbg_0_dbg_uart_0_n_4_3),.ZN(dbg_0_dbg_uart_0_n_4));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b3___05F05d (.D(dbg_0_dbg_uart_0_n_4),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[3]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_49_3 (.A1(dbg_0_dbg_uart_0_n_49_2),.A2(dbg_0_dbg_uart_0_xfer_buf[12]),.B1(dbg_0_dbg_uart_0_n_49_1),.B2(dbg_0_dbg_uart_0_xfer_buf[3]),.ZN(dbg_0_dbg_uart_0_n_49_3));
	INV_X1_LVT dbg_0dbg_uart_0i_49_4 (.A(dbg_0_dbg_uart_0_n_49_3),.ZN(dbg_0_dbg_din[0]));
	INV_X1_LVT dbg_0dbg_uart_0i_52_0 (.A(dbg_0_mem_burst),.ZN(dbg_0_dbg_uart_0_n_52_0));
	INV_X1_LVT dbg_0dbg_uart_0i_50_0 (.A(dbg_0_mem_burst_rd),.ZN(dbg_0_dbg_uart_0_n_50_0));
	INV_X1_LVT dbg_0dbg_uart_0i_50_1 (.A(dbg_0_dbg_uart_0_cmd_valid),.ZN(dbg_0_dbg_uart_0_n_50_1));
	OAI21_X1_LVT dbg_0dbg_uart_0i_50_2 (.A(dbg_0_dbg_uart_0_n_50_0),.B1(dbg_0_dbg_uart_0_n_50_1),.B2(dbg_0_dbg_uart_0_xfer_buf[0]),.ZN(dbg_0_dbg_uart_0_n_132));
	NOR3_X1_LVT dbg_0dbg_uart_0i_13_8 (.A1(dbg_0_dbg_uart_0_n_13_2),.A2(dbg_0_dbg_uart_0_n_13_1),.A3(dbg_0_dbg_uart_0_uart_state[1]),.ZN(dbg_0_dbg_uart_0_n_30));
	AND2_X1_LVT dbg_0dbg_uart_0i_51_0 (.A1(dbg_0_dbg_uart_0_xfer_done),.A2(dbg_0_dbg_uart_0_n_30),.ZN(dbg_0_dbg_uart_0_n_133));
	AOI22_X1_LVT dbg_0dbg_uart_0i_52_1 (.A1(dbg_0_dbg_uart_0_n_52_0),.A2(dbg_0_dbg_uart_0_n_132),.B1(dbg_0_dbg_uart_0_n_133),.B2(dbg_0_mem_burst),.ZN(dbg_0_dbg_uart_0_n_52_1));
	INV_X1_LVT dbg_0dbg_uart_0i_52_2 (.A(dbg_0_dbg_uart_0_n_52_1),.ZN(dbg_0_dbg_rd));
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_4 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[3]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[1]),.ZN(dbg_0_dbg_uart_0_n_4_2));
	INV_X1_LVT dbg_0dbg_uart_0i_4_5 (.A(dbg_0_dbg_uart_0_n_4_2),.ZN(dbg_0_dbg_uart_0_n_3));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b2___05F05d (.D(dbg_0_dbg_uart_0_n_3),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[2]),.QN());
	AOI22_X1_LVT dbg_0dbg_uart_0i_4_2 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[2]),.B1(dbg_0_dbg_rd_rdy),.B2(dbg_0_dbg_dout[0]),.ZN(dbg_0_dbg_uart_0_n_4_1));
	INV_X1_LVT dbg_0dbg_uart_0i_4_3 (.A(dbg_0_dbg_uart_0_n_4_1),.ZN(dbg_0_dbg_uart_0_n_2));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b1___05F05d (.D(dbg_0_dbg_uart_0_n_2),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[1]),.QN());
	AND2_X1_LVT dbg_0dbg_uart_0i_4_1 (.A1(dbg_0_dbg_uart_0_n_4_0),.A2(dbg_0_dbg_uart_0_xfer_buf[1]),.ZN(dbg_0_dbg_uart_0_n_1));
	DFFR_X1_LVT dbg_0dbg_uart_0xfer_buf_reg___05F05b0___05F05d (.D(dbg_0_dbg_uart_0_n_1),.RN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_0),.Q(dbg_0_dbg_uart_0_xfer_buf[0]),.QN());
	OAI21_X1_LVT dbg_0dbg_uart_0i_54_0 (.A(dbg_0_dbg_uart_0_xfer_bit_inc),.B1(dbg_0_dbg_uart_0_n_28),.B2(dbg_0_dbg_uart_0_n_30),.ZN(dbg_0_dbg_uart_0_n_54_0));
	INV_X1_LVT dbg_0dbg_uart_0i_54_1 (.A(dbg_0_dbg_uart_0_n_54_0),.ZN(dbg_0_dbg_uart_0_n_135));
	CLKGATETST_X1_LVT dbg_0dbg_uart_0clk_gate_dbg_uart_txd_reg (.CK(dbg_clk),.E(dbg_0_dbg_uart_0_n_135),.SE(1'b0),.GCK(dbg_0_dbg_uart_0_n_134));
	DFFS_X1_LVT dbg_0dbg_uart_0dbg_uart_txd_reg (.D(dbg_0_dbg_uart_0_xfer_buf[0]),.SN(dbg_0_dbg_uart_0_n_130),.CK(dbg_0_dbg_uart_0_n_134),.Q(dbg_uart_txd),.QN());
	AND2_X1_LVT dbg_0dbg_uart_0i_56_0 (.A1(dbg_0_dbg_uart_0_xfer_done),.A2(dbg_0_dbg_uart_0_n_26),.ZN(dbg_0_dbg_wr));
	CLKGATETST_X1_LVT dbg_0clk_gate_cpu_ctl_reg (.CK(dbg_clk),.E(dbg_0_cpu_ctl_wr),.SE(1'b0),.GCK(dbg_0_n_103));
	DFFR_X1_LVT dbg_0cpu_ctl_reg___05F05b6___05F05d (.D(dbg_0_dbg_din[6]),.RN(dbg_0_n_104),.CK(dbg_0_n_103),.Q(dbg_cpu_reset),.QN());
	INV_X1_LVT dbg_0i_53_0 (.A(cpu_en_s),.ZN(dbg_0_n_53_0));
	OAI21_X1_LVT dbg_0i_53_1 (.A(cpu_halt_st),.B1(dbg_0_n_53_0),.B2(dbg_0_cpu_ctl[1]),.ZN(dbg_0_n_53_1));
	INV_X1_LVT dbg_0i_53_2 (.A(dbg_0_n_53_1),.ZN(dbg_freeze));
	INV_X1_LVT dbg_0i_55_0 (.A(cpu_halt_st),.ZN(dbg_0_n_55_0));
	NAND3_X1_LVT dbg_0i_55_1 (.A1(dbg_0_n_55_0),.A2(dbg_0_cpu_ctl_wr),.A3(dbg_0_dbg_din[0]),.ZN(dbg_0_n_55_1));
	INV_X1_LVT dbg_0i_55_2 (.A(dbg_0_mem_state_nxt_reg[1]),.ZN(dbg_0_n_55_2));
	NOR2_X1_LVT dbg_0i_12_3 (.A1(dbg_0_mem_state[0]),.A2(dbg_0_mem_state[1]),.ZN(dbg_0_n_8));
	NAND3_X1_LVT dbg_0i_55_3 (.A1(dbg_0_n_55_2),.A2(dbg_0_mem_state_nxt_reg[0]),.A3(dbg_0_n_8),.ZN(dbg_0_n_55_3));
	NAND3_X1_LVT dbg_0i_55_4 (.A1(puc_pnd_set),.A2(dbg_0_cpu_ctl[2]),.A3(dbg_en_s),.ZN(dbg_0_n_55_4));
	INV_X1_LVT dbg_0i_55_5 (.A(dbg_0_dbg_swbrk),.ZN(dbg_0_n_55_5));
	NAND4_X1_LVT dbg_0i_55_6 (.A1(dbg_0_n_55_1),.A2(dbg_0_n_55_3),.A3(dbg_0_n_55_4),.A4(dbg_0_n_55_5),.ZN(dbg_0_halt_flag_set));
	INV_X1_LVT dbg_0i_59_0 (.A(dbg_0_halt_flag_set),.ZN(dbg_0_n_59_0));
	INV_X1_LVT dbg_0i_57_0 (.A(dbg_0_n_7),.ZN(dbg_0_n_57_0));
	NOR3_X1_LVT dbg_0i_57_1 (.A1(dbg_0_n_57_0),.A2(dbg_0_mem_state_nxt_reg[0]),.A3(dbg_0_mem_state_nxt_reg[1]),.ZN(dbg_0_n_57_1));
	AND2_X1_LVT dbg_0i_56_0 (.A1(cpu_halt_st),.A2(dbg_0_cpu_ctl_wr),.ZN(dbg_0_n_108));
	AOI21_X1_LVT dbg_0i_57_2 (.A(dbg_0_n_57_1),.B1(dbg_0_dbg_din[1]),.B2(dbg_0_n_108),.ZN(dbg_0_n_57_2));
	INV_X1_LVT dbg_0i_57_3 (.A(dbg_0_n_57_2),.ZN(dbg_0_halt_flag_clr));
	NOR2_X1_LVT dbg_0i_59_1 (.A1(dbg_0_n_59_0),.A2(dbg_0_halt_flag_clr),.ZN(dbg_0_n_110));
	INV_X1_LVT dbg_0i_60_1 (.A(dbg_0_halt_flag_set),.ZN(dbg_0_n_60_1));
	INV_X1_LVT dbg_0i_60_0 (.A(dbg_0_halt_flag_clr),.ZN(dbg_0_n_60_0));
	NAND2_X1_LVT dbg_0i_60_2 (.A1(dbg_0_n_60_1),.A2(dbg_0_n_60_0),.ZN(dbg_0_n_111));
	CLKGATETST_X1_LVT dbg_0clk_gate_halt_flag_reg (.CK(dbg_clk),.E(dbg_0_n_111),.SE(1'b0),.GCK(dbg_0_n_109));
	DFFR_X1_LVT dbg_0halt_flag_reg (.D(dbg_0_n_110),.RN(dbg_0_n_104),.CK(dbg_0_n_109),.Q(dbg_0_halt_flag),.QN());
	NOR2_X1_LVT dbg_0i_66_0 (.A1(dbg_0_halt_flag),.A2(dbg_0_halt_flag_set),.ZN(dbg_0_n_66_0));
	AND2_X1_LVT dbg_0i_62_0 (.A1(dbg_0_dbg_din[2]),.A2(dbg_0_n_108),.ZN(dbg_0_istep));
	DFFR_X1_LVT dbg_0inc_step_reg___05F05b0___05F05d (.D(dbg_0_istep),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_n_113),.QN());
	INV_X1_LVT dbg_0i_64_1 (.A(dbg_0_n_113),.ZN(dbg_0_n_64_1));
	INV_X1_LVT dbg_0i_64_0 (.A(dbg_0_istep),.ZN(dbg_0_n_64_0));
	NAND2_X1_LVT dbg_0i_64_2 (.A1(dbg_0_n_64_1),.A2(dbg_0_n_64_0),.ZN(dbg_0_n_114));
	DFFR_X1_LVT dbg_0inc_step_reg___05F05b1___05F05d (.D(dbg_0_n_114),.RN(dbg_0_n_104),.CK(dbg_clk),.Q(dbg_0_n_112),.QN());
	NOR2_X1_LVT dbg_0i_66_1 (.A1(dbg_0_n_66_0),.A2(dbg_0_n_112),.ZN(dbg_halt_cmd));
	NAND2_X1_LVT dbg_0i_74_18 (.A1(dbg_mem_addr[0]),.A2(dbg_0_mem_ctl[2]),.ZN(dbg_0_n_74_10));
	INV_X1_LVT dbg_0i_74_16 (.A(dbg_0_mem_data[7]),.ZN(dbg_0_n_74_9));
	INV_X1_LVT dbg_0i_74_33 (.A(dbg_0_mem_data[15]),.ZN(dbg_0_n_74_18));
	OAI22_X1_LVT dbg_0i_74_34 (.A1(dbg_0_n_74_10),.A2(dbg_0_n_74_9),.B1(dbg_0_mem_ctl[2]),.B2(dbg_0_n_74_18),.ZN(dbg_mem_dout[15]));
	INV_X1_LVT dbg_0i_74_14 (.A(dbg_0_mem_data[6]),.ZN(dbg_0_n_74_8));
	INV_X1_LVT dbg_0i_74_31 (.A(dbg_0_mem_data[14]),.ZN(dbg_0_n_74_17));
	OAI22_X1_LVT dbg_0i_74_32 (.A1(dbg_0_n_74_10),.A2(dbg_0_n_74_8),.B1(dbg_0_mem_ctl[2]),.B2(dbg_0_n_74_17),.ZN(dbg_mem_dout[14]));
	INV_X1_LVT dbg_0i_74_12 (.A(dbg_0_mem_data[5]),.ZN(dbg_0_n_74_7));
	INV_X1_LVT dbg_0i_74_29 (.A(dbg_0_mem_data[13]),.ZN(dbg_0_n_74_16));
	OAI22_X1_LVT dbg_0i_74_30 (.A1(dbg_0_n_74_10),.A2(dbg_0_n_74_7),.B1(dbg_0_mem_ctl[2]),.B2(dbg_0_n_74_16),.ZN(dbg_mem_dout[13]));
	INV_X1_LVT dbg_0i_74_10 (.A(dbg_0_mem_data[4]),.ZN(dbg_0_n_74_6));
	INV_X1_LVT dbg_0i_74_27 (.A(dbg_0_mem_data[12]),.ZN(dbg_0_n_74_15));
	OAI22_X1_LVT dbg_0i_74_28 (.A1(dbg_0_n_74_10),.A2(dbg_0_n_74_6),.B1(dbg_0_mem_ctl[2]),.B2(dbg_0_n_74_15),.ZN(dbg_mem_dout[12]));
	INV_X1_LVT dbg_0i_74_8 (.A(dbg_0_mem_data[3]),.ZN(dbg_0_n_74_5));
	INV_X1_LVT dbg_0i_74_25 (.A(dbg_0_mem_data[11]),.ZN(dbg_0_n_74_14));
	OAI22_X1_LVT dbg_0i_74_26 (.A1(dbg_0_n_74_10),.A2(dbg_0_n_74_5),.B1(dbg_0_mem_ctl[2]),.B2(dbg_0_n_74_14),.ZN(dbg_mem_dout[11]));
	INV_X1_LVT dbg_0i_74_6 (.A(dbg_0_mem_data[2]),.ZN(dbg_0_n_74_4));
	INV_X1_LVT dbg_0i_74_23 (.A(dbg_0_mem_data[10]),.ZN(dbg_0_n_74_13));
	OAI22_X1_LVT dbg_0i_74_24 (.A1(dbg_0_n_74_10),.A2(dbg_0_n_74_4),.B1(dbg_0_mem_ctl[2]),.B2(dbg_0_n_74_13),.ZN(dbg_mem_dout[10]));
	INV_X1_LVT dbg_0i_74_4 (.A(dbg_0_mem_data[1]),.ZN(dbg_0_n_74_3));
	INV_X1_LVT dbg_0i_74_21 (.A(dbg_0_mem_data[9]),.ZN(dbg_0_n_74_12));
	OAI22_X1_LVT dbg_0i_74_22 (.A1(dbg_0_n_74_10),.A2(dbg_0_n_74_3),.B1(dbg_0_mem_ctl[2]),.B2(dbg_0_n_74_12),.ZN(dbg_mem_dout[9]));
	INV_X1_LVT dbg_0i_74_2 (.A(dbg_0_mem_data[0]),.ZN(dbg_0_n_74_2));
	INV_X1_LVT dbg_0i_74_19 (.A(dbg_0_mem_data[8]),.ZN(dbg_0_n_74_11));
	OAI22_X1_LVT dbg_0i_74_20 (.A1(dbg_0_n_74_10),.A2(dbg_0_n_74_2),.B1(dbg_0_mem_ctl[2]),.B2(dbg_0_n_74_11),.ZN(dbg_mem_dout[8]));
	INV_X1_LVT dbg_0i_74_1 (.A(dbg_mem_addr[0]),.ZN(dbg_0_n_74_1));
	INV_X1_LVT dbg_0i_74_0 (.A(dbg_0_mem_ctl[2]),.ZN(dbg_0_n_74_0));
	NOR2_X1_LVT dbg_0i_74_35 (.A1(dbg_0_n_74_1),.A2(dbg_0_n_74_0),.ZN(dbg_0_n_74_19));
	NOR2_X1_LVT dbg_0i_74_17 (.A1(dbg_0_n_74_19),.A2(dbg_0_n_74_9),.ZN(dbg_mem_dout[7]));
	NOR2_X1_LVT dbg_0i_74_15 (.A1(dbg_0_n_74_19),.A2(dbg_0_n_74_8),.ZN(dbg_mem_dout[6]));
	NOR2_X1_LVT dbg_0i_74_13 (.A1(dbg_0_n_74_19),.A2(dbg_0_n_74_7),.ZN(dbg_mem_dout[5]));
	NOR2_X1_LVT dbg_0i_74_11 (.A1(dbg_0_n_74_19),.A2(dbg_0_n_74_6),.ZN(dbg_mem_dout[4]));
	NOR2_X1_LVT dbg_0i_74_9 (.A1(dbg_0_n_74_19),.A2(dbg_0_n_74_5),.ZN(dbg_mem_dout[3]));
	NOR2_X1_LVT dbg_0i_74_7 (.A1(dbg_0_n_74_19),.A2(dbg_0_n_74_4),.ZN(dbg_mem_dout[2]));
	NOR2_X1_LVT dbg_0i_74_5 (.A1(dbg_0_n_74_19),.A2(dbg_0_n_74_3),.ZN(dbg_mem_dout[1]));
	NOR2_X1_LVT dbg_0i_74_3 (.A1(dbg_0_n_74_19),.A2(dbg_0_n_74_2),.ZN(dbg_mem_dout[0]));
	OR2_X1_LVT multiplier_0i_5_0 (.A1(per_we[0]),.A2(per_we[1]),.ZN(multiplier_0_n_15));
	NAND4_X1_LVT multiplier_0i_0_0 (.A1(per_addr[3]),.A2(per_addr[4]),.A3(per_addr[7]),.A4(per_en),.ZN(multiplier_0_n_0_0));
	NOR4_X1_LVT multiplier_0i_0_1 (.A1(multiplier_0_n_0_0),.A2(per_addr[11]),.A3(per_addr[12]),.A4(per_addr[13]),.ZN(multiplier_0_n_0_1));
	NOR4_X1_LVT multiplier_0i_0_2 (.A1(per_addr[6]),.A2(per_addr[8]),.A3(per_addr[9]),.A4(per_addr[10]),.ZN(multiplier_0_n_0_2));
	NAND2_X1_LVT multiplier_0i_0_3 (.A1(multiplier_0_n_0_1),.A2(multiplier_0_n_0_2),.ZN(multiplier_0_n_0_3));
	NOR2_X1_LVT multiplier_0i_0_4 (.A1(multiplier_0_n_0_3),.A2(per_addr[5]),.ZN(multiplier_0_reg_sel));
	AND2_X1_LVT multiplier_0i_6_0 (.A1(multiplier_0_n_15),.A2(multiplier_0_reg_sel),.ZN(multiplier_0_reg_write));
	INV_X1_LVT multiplier_0i_3_6 (.A(per_addr[2]),.ZN(multiplier_0_n_3_2));
	NOR3_X1_LVT multiplier_0i_3_7 (.A1(multiplier_0_n_3_2),.A2(per_addr[0]),.A3(per_addr[1]),.ZN(multiplier_0_n_5));
	AND2_X1_LVT multiplier_0i_7_4 (.A1(multiplier_0_reg_write),.A2(multiplier_0_n_5),.ZN(multiplier_0_op2_wr));
	INV_X1_LVT multiplier_0i_21_0 (.A(puc_rst),.ZN(multiplier_0_n_38));
	DFFR_X1_LVT multiplier_0cycle_reg___05F05b0___05F05d (.D(multiplier_0_op2_wr),.RN(multiplier_0_n_38),.CK(mclk),.Q(multiplier_0_cycle[0]),.QN());
	DFFR_X1_LVT multiplier_0cycle_reg___05F05b1___05F05d (.D(multiplier_0_cycle[0]),.RN(multiplier_0_n_38),.CK(mclk),.Q(multiplier_0_cycle[1]),.QN());
	INV_X1_LVT multiplier_0i_60_0 (.A(multiplier_0_cycle[1]),.ZN(multiplier_0_n_60_0));
	INV_X1_LVT multiplier_0i_38_0 (.A(multiplier_0_op2_wr),.ZN(multiplier_0_n_38_0));
	INV_X1_LVT multiplier_0i_3_3 (.A(per_addr[1]),.ZN(multiplier_0_n_3_1));
	NOR3_X1_LVT multiplier_0i_3_4 (.A1(multiplier_0_n_3_1),.A2(per_addr[0]),.A3(per_addr[2]),.ZN(multiplier_0_n_3));
	AND2_X1_LVT multiplier_0i_7_2 (.A1(multiplier_0_reg_write),.A2(multiplier_0_n_3),.ZN(multiplier_0_n_18));
	INV_X1_LVT multiplier_0i_3_1 (.A(per_addr[0]),.ZN(multiplier_0_n_3_0));
	NOR3_X1_LVT multiplier_0i_3_5 (.A1(multiplier_0_n_3_1),.A2(multiplier_0_n_3_0),.A3(per_addr[2]),.ZN(multiplier_0_n_4));
	AND2_X1_LVT multiplier_0i_7_3 (.A1(multiplier_0_reg_write),.A2(multiplier_0_n_4),.ZN(multiplier_0_n_19));
	OR2_X1_LVT multiplier_0i_36_0 (.A1(multiplier_0_n_18),.A2(multiplier_0_n_19),.ZN(multiplier_0_n_68));
	NOR3_X1_LVT multiplier_0i_3_0 (.A1(per_addr[0]),.A2(per_addr[1]),.A3(per_addr[2]),.ZN(multiplier_0_n_1));
	AND2_X1_LVT multiplier_0i_7_0 (.A1(multiplier_0_n_1),.A2(multiplier_0_reg_write),.ZN(multiplier_0_n_16));
	NOR3_X1_LVT multiplier_0i_3_2 (.A1(multiplier_0_n_3_0),.A2(per_addr[1]),.A3(per_addr[2]),.ZN(multiplier_0_n_2));
	AND2_X1_LVT multiplier_0i_7_1 (.A1(multiplier_0_reg_write),.A2(multiplier_0_n_2),.ZN(multiplier_0_n_17));
	OR4_X1_LVT multiplier_0i_24_0 (.A1(multiplier_0_n_16),.A2(multiplier_0_n_19),.A3(multiplier_0_n_18),.A4(multiplier_0_n_17),.ZN(multiplier_0_op1_wr));
	CLKGATETST_X1_LVT multiplier_0clk_gate_acc_sel_reg (.CK(mclk),.E(multiplier_0_op1_wr),.SE(1'b0),.GCK(multiplier_0_n_67));
	DFFR_X1_LVT multiplier_0acc_sel_reg (.D(multiplier_0_n_68),.RN(multiplier_0_n_38),.CK(multiplier_0_n_67),.Q(multiplier_0_acc_sel),.QN());
	NOR2_X1_LVT multiplier_0i_38_1 (.A1(multiplier_0_n_38_0),.A2(multiplier_0_acc_sel),.ZN(multiplier_0_result_clr));
	NOR3_X1_LVT multiplier_0i_3_8 (.A1(multiplier_0_n_3_2),.A2(multiplier_0_n_3_0),.A3(per_addr[1]),.ZN(multiplier_0_n_6));
	AND2_X1_LVT multiplier_0i_7_5 (.A1(multiplier_0_reg_write),.A2(multiplier_0_n_6),.ZN(multiplier_0_reslo_wr));
	NOR2_X1_LVT multiplier_0i_45_0 (.A1(multiplier_0_result_clr),.A2(multiplier_0_reslo_wr),.ZN(multiplier_0_n_45_0));
	INV_X1_LVT multiplier_0i_34_16 (.A(multiplier_0_cycle[0]),.ZN(multiplier_0_n_34_8));
	INV_X1_LVT multiplier_0i_29_0 (.A(multiplier_0_cycle[0]),.ZN(multiplier_0_n_29_0));
	CLKGATETST_X1_LVT multiplier_0clk_gate_op2_reg (.CK(mclk),.E(multiplier_0_op2_wr),.SE(1'b0),.GCK(multiplier_0_n_20));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b4___05F05d (.D(per_din[4]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_20),.Q(multiplier_0_op2_reg[4]),.QN());
	AND2_X1_LVT multiplier_0i_8_4 (.A1(per_we[1]),.A2(per_din[12]),.ZN(multiplier_0_per_din_msk[12]));
	CLKGATETST_X1_LVT multiplier_0clk_gate_op2_reg___05F_05F0 (.CK(mclk),.E(multiplier_0_op2_wr),.SE(1'b0),.GCK(multiplier_0_n_21));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b12___05F05d (.D(multiplier_0_per_din_msk[12]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_21),.Q(multiplier_0_op2_reg[12]),.QN());
	AOI22_X1_LVT multiplier_0i_29_9 (.A1(multiplier_0_n_29_0),.A2(multiplier_0_op2_reg[4]),.B1(multiplier_0_cycle[0]),.B2(multiplier_0_op2_reg[12]),.ZN(multiplier_0_n_29_5));
	INV_X1_LVT multiplier_0i_29_10 (.A(multiplier_0_n_29_5),.ZN(multiplier_0_op2_xp[4]));
	CLKGATETST_X1_LVT multiplier_0clk_gate_op1_reg (.CK(mclk),.E(multiplier_0_op1_wr),.SE(1'b0),.GCK(multiplier_0_n_41));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b3___05F05d (.D(per_din[3]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[3]),.QN());
	NAND2_X1_LVT multiplier_0i_32_71 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_32_71));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b3___05F05d (.D(per_din[3]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_20),.Q(multiplier_0_op2_reg[3]),.QN());
	AND2_X1_LVT multiplier_0i_8_3 (.A1(per_we[1]),.A2(per_din[11]),.ZN(multiplier_0_per_din_msk[11]));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b11___05F05d (.D(multiplier_0_per_din_msk[11]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_21),.Q(multiplier_0_op2_reg[11]),.QN());
	AOI22_X1_LVT multiplier_0i_29_7 (.A1(multiplier_0_n_29_0),.A2(multiplier_0_op2_reg[3]),.B1(multiplier_0_cycle[0]),.B2(multiplier_0_op2_reg[11]),.ZN(multiplier_0_n_29_4));
	INV_X1_LVT multiplier_0i_29_8 (.A(multiplier_0_n_29_4),.ZN(multiplier_0_op2_xp[3]));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b4___05F05d (.D(per_din[4]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[4]),.QN());
	NAND2_X1_LVT multiplier_0i_32_55 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_32_55));
	XNOR2_X1_LVT multiplier_0i_32_229 (.A(multiplier_0_n_32_71),.B(multiplier_0_n_32_55),.ZN(multiplier_0_n_32_234));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b2___05F05d (.D(per_din[2]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_20),.Q(multiplier_0_op2_reg[2]),.QN());
	AND2_X1_LVT multiplier_0i_8_2 (.A1(per_we[1]),.A2(per_din[10]),.ZN(multiplier_0_per_din_msk[10]));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b10___05F05d (.D(multiplier_0_per_din_msk[10]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_21),.Q(multiplier_0_op2_reg[10]),.QN());
	AOI22_X1_LVT multiplier_0i_29_5 (.A1(multiplier_0_n_29_0),.A2(multiplier_0_op2_reg[2]),.B1(multiplier_0_cycle[0]),.B2(multiplier_0_op2_reg[10]),.ZN(multiplier_0_n_29_3));
	INV_X1_LVT multiplier_0i_29_6 (.A(multiplier_0_n_29_3),.ZN(multiplier_0_op2_xp[2]));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b5___05F05d (.D(per_din[5]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[5]),.QN());
	NAND2_X1_LVT multiplier_0i_32_39 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_32_39));
	XNOR2_X1_LVT multiplier_0i_32_230 (.A(multiplier_0_n_32_234),.B(multiplier_0_n_32_39),.ZN(multiplier_0_n_32_235));
	INV_X1_LVT multiplier_0i_32_231 (.A(multiplier_0_n_32_235),.ZN(multiplier_0_n_32_236));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b7___05F05d (.D(per_din[7]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_20),.Q(multiplier_0_op2_reg[7]),.QN());
	AND2_X1_LVT multiplier_0i_8_7 (.A1(per_we[1]),.A2(per_din[15]),.ZN(multiplier_0_per_din_msk[15]));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b15___05F05d (.D(multiplier_0_per_din_msk[15]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_21),.Q(multiplier_0_op2_reg[15]),.QN());
	AOI22_X1_LVT multiplier_0i_29_15 (.A1(multiplier_0_n_29_0),.A2(multiplier_0_op2_reg[7]),.B1(multiplier_0_cycle[0]),.B2(multiplier_0_op2_reg[15]),.ZN(multiplier_0_n_29_8));
	INV_X1_LVT multiplier_0i_29_16 (.A(multiplier_0_n_29_8),.ZN(multiplier_0_op2_xp[7]));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b0___05F05d (.D(per_din[0]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[0]),.QN());
	NAND2_X1_LVT multiplier_0i_32_119 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[0]),.ZN(multiplier_0_n_32_119));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b6___05F05d (.D(per_din[6]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_20),.Q(multiplier_0_op2_reg[6]),.QN());
	AND2_X1_LVT multiplier_0i_8_6 (.A1(per_we[1]),.A2(per_din[14]),.ZN(multiplier_0_per_din_msk[14]));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b14___05F05d (.D(multiplier_0_per_din_msk[14]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_21),.Q(multiplier_0_op2_reg[14]),.QN());
	AOI22_X1_LVT multiplier_0i_29_13 (.A1(multiplier_0_n_29_0),.A2(multiplier_0_op2_reg[6]),.B1(multiplier_0_cycle[0]),.B2(multiplier_0_op2_reg[14]),.ZN(multiplier_0_n_29_7));
	INV_X1_LVT multiplier_0i_29_14 (.A(multiplier_0_n_29_7),.ZN(multiplier_0_op2_xp[6]));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b1___05F05d (.D(per_din[1]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[1]),.QN());
	NAND2_X1_LVT multiplier_0i_32_103 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_32_103));
	XNOR2_X1_LVT multiplier_0i_32_222 (.A(multiplier_0_n_32_119),.B(multiplier_0_n_32_103),.ZN(multiplier_0_n_32_227));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b5___05F05d (.D(per_din[5]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_20),.Q(multiplier_0_op2_reg[5]),.QN());
	AND2_X1_LVT multiplier_0i_8_5 (.A1(per_we[1]),.A2(per_din[13]),.ZN(multiplier_0_per_din_msk[13]));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b13___05F05d (.D(multiplier_0_per_din_msk[13]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_21),.Q(multiplier_0_op2_reg[13]),.QN());
	AOI22_X1_LVT multiplier_0i_29_11 (.A1(multiplier_0_n_29_0),.A2(multiplier_0_op2_reg[5]),.B1(multiplier_0_cycle[0]),.B2(multiplier_0_op2_reg[13]),.ZN(multiplier_0_n_29_6));
	INV_X1_LVT multiplier_0i_29_12 (.A(multiplier_0_n_29_6),.ZN(multiplier_0_op2_xp[5]));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b2___05F05d (.D(per_din[2]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[2]),.QN());
	NAND2_X1_LVT multiplier_0i_32_87 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_32_87));
	XNOR2_X1_LVT multiplier_0i_32_223 (.A(multiplier_0_n_32_227),.B(multiplier_0_n_32_87),.ZN(multiplier_0_n_32_228));
	INV_X1_LVT multiplier_0i_32_224 (.A(multiplier_0_n_32_228),.ZN(multiplier_0_n_32_229));
	NAND2_X1_LVT multiplier_0i_32_85 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[0]),.ZN(multiplier_0_n_32_85));
	NAND2_X1_LVT multiplier_0i_32_69 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_32_69));
	XNOR2_X1_LVT multiplier_0i_32_182 (.A(multiplier_0_n_32_85),.B(multiplier_0_n_32_69),.ZN(multiplier_0_n_32_183));
	NAND2_X1_LVT multiplier_0i_32_53 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_32_53));
	XNOR2_X1_LVT multiplier_0i_32_183 (.A(multiplier_0_n_32_183),.B(multiplier_0_n_32_53),.ZN(multiplier_0_n_32_184));
	INV_X1_LVT multiplier_0i_32_184 (.A(multiplier_0_n_32_184),.ZN(multiplier_0_n_32_185));
	NAND2_X1_LVT multiplier_0i_32_35 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_32_35));
	NAND2_X1_LVT multiplier_0i_32_51 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[0]),.ZN(multiplier_0_n_32_51));
	NOR2_X1_LVT multiplier_0i_32_159 (.A1(multiplier_0_n_32_35),.A2(multiplier_0_n_32_51),.ZN(multiplier_0_n_32_159));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b1___05F05d (.D(per_din[1]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_20),.Q(multiplier_0_op2_reg[1]),.QN());
	AND2_X1_LVT multiplier_0i_8_1 (.A1(per_we[1]),.A2(per_din[9]),.ZN(multiplier_0_per_din_msk[9]));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b9___05F05d (.D(multiplier_0_per_din_msk[9]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_21),.Q(multiplier_0_op2_reg[9]),.QN());
	AOI22_X1_LVT multiplier_0i_29_3 (.A1(multiplier_0_n_29_0),.A2(multiplier_0_op2_reg[1]),.B1(multiplier_0_cycle[0]),.B2(multiplier_0_op2_reg[9]),.ZN(multiplier_0_n_29_2));
	INV_X1_LVT multiplier_0i_29_4 (.A(multiplier_0_n_29_2),.ZN(multiplier_0_op2_xp[1]));
	NAND2_X1_LVT multiplier_0i_32_19 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_32_19));
	NOR2_X1_LVT multiplier_0i_32_160 (.A1(multiplier_0_n_32_19),.A2(multiplier_0_n_32_51),.ZN(multiplier_0_n_32_160));
	NOR2_X1_LVT multiplier_0i_32_161 (.A1(multiplier_0_n_32_19),.A2(multiplier_0_n_32_35),.ZN(multiplier_0_n_32_161));
	OR3_X1_LVT multiplier_0i_32_158 (.A1(multiplier_0_n_32_159),.A2(multiplier_0_n_32_160),.A3(multiplier_0_n_32_161),.ZN(multiplier_0_n_32_158));
	NAND2_X1_LVT multiplier_0i_32_20 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_32_20));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b0___05F05d (.D(per_din[0]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_20),.Q(multiplier_0_op2_reg[0]),.QN());
	AND2_X1_LVT multiplier_0i_8_0 (.A1(per_din[8]),.A2(per_we[1]),.ZN(multiplier_0_per_din_msk[8]));
	DFFR_X1_LVT multiplier_0op2_reg___05F05b8___05F05d (.D(multiplier_0_per_din_msk[8]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_21),.Q(multiplier_0_op2_reg[8]),.QN());
	AOI22_X1_LVT multiplier_0i_29_1 (.A1(multiplier_0_n_29_0),.A2(multiplier_0_op2_reg[0]),.B1(multiplier_0_op2_reg[8]),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_n_29_1));
	INV_X1_LVT multiplier_0i_29_2 (.A(multiplier_0_n_29_1),.ZN(multiplier_0_op2_xp[0]));
	NAND2_X1_LVT multiplier_0i_32_4 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_32_4));
	XNOR2_X1_LVT multiplier_0i_32_173 (.A(multiplier_0_n_32_20),.B(multiplier_0_n_32_4),.ZN(multiplier_0_n_32_173));
	NAND2_X1_LVT multiplier_0i_32_18 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_32_18));
	NAND2_X1_LVT multiplier_0i_32_34 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[0]),.ZN(multiplier_0_n_32_34));
	NOR2_X1_LVT multiplier_0i_32_154 (.A1(multiplier_0_n_32_18),.A2(multiplier_0_n_32_34),.ZN(multiplier_0_n_32_154));
	NAND2_X1_LVT multiplier_0i_32_3 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_32_3));
	INV_X1_LVT multiplier_0i_32_164 (.A(multiplier_0_n_32_3),.ZN(multiplier_0_n_32_164));
	NAND2_X1_LVT multiplier_0i_32_163 (.A1(multiplier_0_n_32_154),.A2(multiplier_0_n_32_164),.ZN(multiplier_0_n_32_163));
	INV_X1_LVT multiplier_0i_32_165 (.A(multiplier_0_n_32_163),.ZN(multiplier_0_n_32_165));
	XNOR2_X1_LVT multiplier_0i_32_174 (.A(multiplier_0_n_32_173),.B(multiplier_0_n_32_165),.ZN(multiplier_0_n_32_174));
	HA_X1_LVT multiplier_0i_32_181 (.A(multiplier_0_n_32_158),.B(multiplier_0_n_32_174),.CO(multiplier_0_n_32_182),.S(multiplier_0_n_32_181));
	HA_X1_LVT multiplier_0i_32_197 (.A(multiplier_0_n_32_185),.B(multiplier_0_n_32_182),.CO(multiplier_0_n_32_200),.S(multiplier_0_n_32_199));
	NAND2_X1_LVT multiplier_0i_32_52 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_32_52));
	NAND2_X1_LVT multiplier_0i_32_68 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[0]),.ZN(multiplier_0_n_32_68));
	NOR2_X1_LVT multiplier_0i_32_170 (.A1(multiplier_0_n_32_52),.A2(multiplier_0_n_32_68),.ZN(multiplier_0_n_32_170));
	NAND2_X1_LVT multiplier_0i_32_36 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_32_36));
	NOR2_X1_LVT multiplier_0i_32_171 (.A1(multiplier_0_n_32_36),.A2(multiplier_0_n_32_68),.ZN(multiplier_0_n_32_171));
	NOR2_X1_LVT multiplier_0i_32_172 (.A1(multiplier_0_n_32_36),.A2(multiplier_0_n_32_52),.ZN(multiplier_0_n_32_172));
	OR3_X1_LVT multiplier_0i_32_169 (.A1(multiplier_0_n_32_170),.A2(multiplier_0_n_32_171),.A3(multiplier_0_n_32_172),.ZN(multiplier_0_n_32_169));
	OR2_X1_LVT multiplier_0i_32_176 (.A1(multiplier_0_n_32_4),.A2(multiplier_0_n_32_20),.ZN(multiplier_0_n_32_176));
	INV_X1_LVT multiplier_0i_32_178 (.A(multiplier_0_n_32_20),.ZN(multiplier_0_n_32_178));
	NAND2_X1_LVT multiplier_0i_32_177 (.A1(multiplier_0_n_32_165),.A2(multiplier_0_n_32_178),.ZN(multiplier_0_n_32_177));
	INV_X1_LVT multiplier_0i_32_180 (.A(multiplier_0_n_32_4),.ZN(multiplier_0_n_32_180));
	NAND2_X1_LVT multiplier_0i_32_179 (.A1(multiplier_0_n_32_165),.A2(multiplier_0_n_32_180),.ZN(multiplier_0_n_32_179));
	NAND3_X1_LVT multiplier_0i_32_175 (.A1(multiplier_0_n_32_176),.A2(multiplier_0_n_32_177),.A3(multiplier_0_n_32_179),.ZN(multiplier_0_n_32_175));
	NAND2_X1_LVT multiplier_0i_32_37 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_32_37));
	NAND2_X1_LVT multiplier_0i_32_21 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_32_21));
	XNOR2_X1_LVT multiplier_0i_32_189 (.A(multiplier_0_n_32_37),.B(multiplier_0_n_32_21),.ZN(multiplier_0_n_32_190));
	NAND2_X1_LVT multiplier_0i_32_5 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_32_5));
	XNOR2_X1_LVT multiplier_0i_32_190 (.A(multiplier_0_n_32_190),.B(multiplier_0_n_32_5),.ZN(multiplier_0_n_32_191));
	INV_X1_LVT multiplier_0i_32_191 (.A(multiplier_0_n_32_191),.ZN(multiplier_0_n_32_192));
	FA_X1_LVT multiplier_0i_32_196 (.A(multiplier_0_n_32_169),.B(multiplier_0_n_32_175),.CI(multiplier_0_n_32_192),.CO(multiplier_0_n_32_198),.S(multiplier_0_n_32_197));
	HA_X1_LVT multiplier_0i_32_221 (.A(multiplier_0_n_32_200),.B(multiplier_0_n_32_198),.CO(multiplier_0_n_32_226),.S(multiplier_0_n_32_225));
	FA_X1_LVT multiplier_0i_32_245 (.A(multiplier_0_n_32_236),.B(multiplier_0_n_32_229),.CI(multiplier_0_n_32_226),.CO(multiplier_0_n_32_252),.S(multiplier_0_n_32_251));
	NAND2_X1_LVT multiplier_0i_32_86 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_32_86));
	NAND2_X1_LVT multiplier_0i_32_102 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[0]),.ZN(multiplier_0_n_32_102));
	NOR2_X1_LVT multiplier_0i_32_202 (.A1(multiplier_0_n_32_86),.A2(multiplier_0_n_32_102),.ZN(multiplier_0_n_32_205));
	NAND2_X1_LVT multiplier_0i_32_70 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_32_70));
	NOR2_X1_LVT multiplier_0i_32_203 (.A1(multiplier_0_n_32_70),.A2(multiplier_0_n_32_102),.ZN(multiplier_0_n_32_206));
	NOR2_X1_LVT multiplier_0i_32_204 (.A1(multiplier_0_n_32_70),.A2(multiplier_0_n_32_86),.ZN(multiplier_0_n_32_207));
	OR3_X1_LVT multiplier_0i_32_201 (.A1(multiplier_0_n_32_205),.A2(multiplier_0_n_32_206),.A3(multiplier_0_n_32_207),.ZN(multiplier_0_n_32_204));
	NOR2_X1_LVT multiplier_0i_32_193 (.A1(multiplier_0_n_32_21),.A2(multiplier_0_n_32_37),.ZN(multiplier_0_n_32_194));
	NOR2_X1_LVT multiplier_0i_32_194 (.A1(multiplier_0_n_32_5),.A2(multiplier_0_n_32_37),.ZN(multiplier_0_n_32_195));
	NOR2_X1_LVT multiplier_0i_32_195 (.A1(multiplier_0_n_32_5),.A2(multiplier_0_n_32_21),.ZN(multiplier_0_n_32_196));
	OR3_X1_LVT multiplier_0i_32_192 (.A1(multiplier_0_n_32_194),.A2(multiplier_0_n_32_195),.A3(multiplier_0_n_32_196),.ZN(multiplier_0_n_32_193));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b6___05F05d (.D(per_din[6]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[6]),.QN());
	NAND2_X1_LVT multiplier_0i_32_6 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_32_6));
	INV_X1_LVT multiplier_0i_32_217 (.A(multiplier_0_n_32_6),.ZN(multiplier_0_n_32_220));
	NAND2_X1_LVT multiplier_0i_32_216 (.A1(multiplier_0_n_32_193),.A2(multiplier_0_n_32_220),.ZN(multiplier_0_n_32_219));
	NOR2_X1_LVT multiplier_0i_32_186 (.A1(multiplier_0_n_32_69),.A2(multiplier_0_n_32_85),.ZN(multiplier_0_n_32_187));
	NOR2_X1_LVT multiplier_0i_32_187 (.A1(multiplier_0_n_32_53),.A2(multiplier_0_n_32_85),.ZN(multiplier_0_n_32_188));
	NOR2_X1_LVT multiplier_0i_32_188 (.A1(multiplier_0_n_32_53),.A2(multiplier_0_n_32_69),.ZN(multiplier_0_n_32_189));
	OR3_X1_LVT multiplier_0i_32_185 (.A1(multiplier_0_n_32_187),.A2(multiplier_0_n_32_188),.A3(multiplier_0_n_32_189),.ZN(multiplier_0_n_32_186));
	NAND2_X1_LVT multiplier_0i_32_218 (.A1(multiplier_0_n_32_186),.A2(multiplier_0_n_32_220),.ZN(multiplier_0_n_32_221));
	NAND2_X1_LVT multiplier_0i_32_219 (.A1(multiplier_0_n_32_186),.A2(multiplier_0_n_32_193),.ZN(multiplier_0_n_32_222));
	NAND3_X1_LVT multiplier_0i_32_215 (.A1(multiplier_0_n_32_219),.A2(multiplier_0_n_32_221),.A3(multiplier_0_n_32_222),.ZN(multiplier_0_n_32_218));
	NAND2_X1_LVT multiplier_0i_32_23 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_32_23));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b7___05F05d (.D(per_din[7]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[7]),.QN());
	NAND2_X1_LVT multiplier_0i_32_7 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_32_7));
	XNOR2_X1_LVT multiplier_0i_32_236 (.A(multiplier_0_n_32_23),.B(multiplier_0_n_32_7),.ZN(multiplier_0_n_32_241));
	NAND2_X1_LVT multiplier_0i_32_38 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_32_38));
	NAND2_X1_LVT multiplier_0i_32_54 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_32_54));
	NOR2_X1_LVT multiplier_0i_32_209 (.A1(multiplier_0_n_32_38),.A2(multiplier_0_n_32_54),.ZN(multiplier_0_n_32_212));
	NAND2_X1_LVT multiplier_0i_32_22 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_32_22));
	NOR2_X1_LVT multiplier_0i_32_210 (.A1(multiplier_0_n_32_22),.A2(multiplier_0_n_32_54),.ZN(multiplier_0_n_32_213));
	NOR2_X1_LVT multiplier_0i_32_211 (.A1(multiplier_0_n_32_22),.A2(multiplier_0_n_32_38),.ZN(multiplier_0_n_32_214));
	OR3_X1_LVT multiplier_0i_32_208 (.A1(multiplier_0_n_32_212),.A2(multiplier_0_n_32_213),.A3(multiplier_0_n_32_214),.ZN(multiplier_0_n_32_211));
	XNOR2_X1_LVT multiplier_0i_32_237 (.A(multiplier_0_n_32_241),.B(multiplier_0_n_32_211),.ZN(multiplier_0_n_32_242));
	FA_X1_LVT multiplier_0i_32_244 (.A(multiplier_0_n_32_204),.B(multiplier_0_n_32_218),.CI(multiplier_0_n_32_242),.CO(multiplier_0_n_32_250),.S(multiplier_0_n_32_249));
	XNOR2_X1_LVT multiplier_0i_32_205 (.A(multiplier_0_n_32_54),.B(multiplier_0_n_32_38),.ZN(multiplier_0_n_32_208));
	XNOR2_X1_LVT multiplier_0i_32_206 (.A(multiplier_0_n_32_208),.B(multiplier_0_n_32_22),.ZN(multiplier_0_n_32_209));
	INV_X1_LVT multiplier_0i_32_207 (.A(multiplier_0_n_32_209),.ZN(multiplier_0_n_32_210));
	XNOR2_X1_LVT multiplier_0i_32_198 (.A(multiplier_0_n_32_102),.B(multiplier_0_n_32_86),.ZN(multiplier_0_n_32_201));
	XNOR2_X1_LVT multiplier_0i_32_199 (.A(multiplier_0_n_32_201),.B(multiplier_0_n_32_70),.ZN(multiplier_0_n_32_202));
	INV_X1_LVT multiplier_0i_32_200 (.A(multiplier_0_n_32_202),.ZN(multiplier_0_n_32_203));
	XNOR2_X1_LVT multiplier_0i_32_212 (.A(multiplier_0_n_32_6),.B(multiplier_0_n_32_193),.ZN(multiplier_0_n_32_215));
	XNOR2_X1_LVT multiplier_0i_32_213 (.A(multiplier_0_n_32_215),.B(multiplier_0_n_32_186),.ZN(multiplier_0_n_32_216));
	INV_X1_LVT multiplier_0i_32_214 (.A(multiplier_0_n_32_216),.ZN(multiplier_0_n_32_217));
	FA_X1_LVT multiplier_0i_32_220 (.A(multiplier_0_n_32_210),.B(multiplier_0_n_32_203),.CI(multiplier_0_n_32_217),.CO(multiplier_0_n_32_224),.S(multiplier_0_n_32_223));
	HA_X1_LVT multiplier_0i_32_246 (.A(multiplier_0_n_32_249),.B(multiplier_0_n_32_224),.CO(multiplier_0_n_32_254),.S(multiplier_0_n_32_253));
	XNOR2_X1_LVT multiplier_0i_32_166 (.A(multiplier_0_n_32_68),.B(multiplier_0_n_32_52),.ZN(multiplier_0_n_32_166));
	XNOR2_X1_LVT multiplier_0i_32_167 (.A(multiplier_0_n_32_166),.B(multiplier_0_n_32_36),.ZN(multiplier_0_n_32_167));
	INV_X1_LVT multiplier_0i_32_168 (.A(multiplier_0_n_32_167),.ZN(multiplier_0_n_32_168));
	XNOR2_X1_LVT multiplier_0i_32_162 (.A(multiplier_0_n_32_3),.B(multiplier_0_n_32_154),.ZN(multiplier_0_n_32_162));
	XNOR2_X1_LVT multiplier_0i_32_155 (.A(multiplier_0_n_32_51),.B(multiplier_0_n_32_35),.ZN(multiplier_0_n_32_155));
	XNOR2_X1_LVT multiplier_0i_32_156 (.A(multiplier_0_n_32_155),.B(multiplier_0_n_32_19),.ZN(multiplier_0_n_32_156));
	INV_X1_LVT multiplier_0i_32_157 (.A(multiplier_0_n_32_156),.ZN(multiplier_0_n_32_157));
	XNOR2_X1_LVT multiplier_0i_32_152 (.A(multiplier_0_n_32_34),.B(multiplier_0_n_32_18),.ZN(multiplier_0_n_32_152));
	INV_X1_LVT multiplier_0i_32_153 (.A(multiplier_0_n_32_152),.ZN(multiplier_0_n_32_153));
	NAND2_X1_LVT multiplier_0i_32_2 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_32_2));
	INV_X1_LVT multiplier_0i_32_594 (.A(multiplier_0_n_32_2),.ZN(multiplier_0_n_32_651));
	NAND2_X1_LVT multiplier_0i_32_593 (.A1(multiplier_0_n_32_153),.A2(multiplier_0_n_32_651),.ZN(multiplier_0_n_32_650));
	NAND2_X1_LVT multiplier_0i_32_1 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_32_1));
	NAND2_X1_LVT multiplier_0i_32_17 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[0]),.ZN(multiplier_0_n_32_17));
	NOR2_X1_LVT multiplier_0i_32_588 (.A1(multiplier_0_n_32_1),.A2(multiplier_0_n_32_17),.ZN(multiplier_0_n_32_646));
	NAND2_X1_LVT multiplier_0i_32_595 (.A1(multiplier_0_n_32_646),.A2(multiplier_0_n_32_651),.ZN(multiplier_0_n_32_652));
	NAND2_X1_LVT multiplier_0i_32_596 (.A1(multiplier_0_n_32_646),.A2(multiplier_0_n_32_153),.ZN(multiplier_0_n_32_653));
	NAND3_X1_LVT multiplier_0i_32_592 (.A1(multiplier_0_n_32_650),.A2(multiplier_0_n_32_652),.A3(multiplier_0_n_32_653),.ZN(multiplier_0_n_32_649));
	FA_X1_LVT multiplier_0i_32_597 (.A(multiplier_0_n_32_162),.B(multiplier_0_n_32_157),.CI(multiplier_0_n_32_649),.CO(multiplier_0_n_32_654),.S(multiplier_0_n_45));
	FA_X1_LVT multiplier_0i_32_598 (.A(multiplier_0_n_32_168),.B(multiplier_0_n_32_181),.CI(multiplier_0_n_32_654),.CO(multiplier_0_n_32_655),.S(multiplier_0_n_46));
	FA_X1_LVT multiplier_0i_32_599 (.A(multiplier_0_n_32_197),.B(multiplier_0_n_32_199),.CI(multiplier_0_n_32_655),.CO(multiplier_0_n_32_656),.S(multiplier_0_n_47));
	FA_X1_LVT multiplier_0i_32_600 (.A(multiplier_0_n_32_225),.B(multiplier_0_n_32_223),.CI(multiplier_0_n_32_656),.CO(multiplier_0_n_32_657),.S(multiplier_0_n_48));
	FA_X1_LVT multiplier_0i_32_601 (.A(multiplier_0_n_32_251),.B(multiplier_0_n_32_253),.CI(multiplier_0_n_32_657),.CO(multiplier_0_n_32_658),.S(multiplier_0_n_49));
	INV_X1_LVT multiplier_0i_34_14 (.A(multiplier_0_n_49),.ZN(multiplier_0_n_34_7));
	OR2_X1_LVT multiplier_0i_26_0 (.A1(multiplier_0_n_17),.A2(multiplier_0_n_19),.ZN(multiplier_0_n_40));
	CLKGATETST_X1_LVT multiplier_0clk_gate_sign_sel_reg (.CK(mclk),.E(multiplier_0_op1_wr),.SE(1'b0),.GCK(multiplier_0_n_39));
	DFFR_X1_LVT multiplier_0sign_sel_reg (.D(multiplier_0_n_40),.RN(multiplier_0_n_38),.CK(multiplier_0_n_39),.Q(multiplier_0_sign_sel),.QN());
	AND2_X1_LVT multiplier_0i_28_0 (.A1(multiplier_0_op2_reg[15]),.A2(multiplier_0_sign_sel),.ZN(multiplier_0_op2_hi_xp[8]));
	AND2_X1_LVT multiplier_0i_29_17 (.A1(multiplier_0_cycle[0]),.A2(multiplier_0_op2_hi_xp[8]),.ZN(multiplier_0_op2_xp[8]));
	NAND2_X1_LVT multiplier_0i_32_141 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_32_141));
	NAND2_X1_LVT multiplier_0i_32_125 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_32_125));
	XNOR2_X1_LVT multiplier_0i_32_380 (.A(multiplier_0_n_32_141),.B(multiplier_0_n_32_125),.ZN(multiplier_0_n_32_407));
	NAND2_X1_LVT multiplier_0i_32_109 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_32_109));
	XNOR2_X1_LVT multiplier_0i_32_381 (.A(multiplier_0_n_32_407),.B(multiplier_0_n_32_109),.ZN(multiplier_0_n_32_408));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b11___05F05d (.D(multiplier_0_per_din_msk[11]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[11]),.QN());
	NAND2_X1_LVT multiplier_0i_32_28 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_32_28));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b10___05F05d (.D(multiplier_0_per_din_msk[10]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[10]),.QN());
	NAND2_X1_LVT multiplier_0i_32_44 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_32_44));
	NOR2_X1_LVT multiplier_0i_32_373 (.A1(multiplier_0_n_32_28),.A2(multiplier_0_n_32_44),.ZN(multiplier_0_n_32_396));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b12___05F05d (.D(multiplier_0_per_din_msk[12]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[12]),.QN());
	NAND2_X1_LVT multiplier_0i_32_12 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_32_12));
	NOR2_X1_LVT multiplier_0i_32_374 (.A1(multiplier_0_n_32_12),.A2(multiplier_0_n_32_44),.ZN(multiplier_0_n_32_397));
	NOR2_X1_LVT multiplier_0i_32_375 (.A1(multiplier_0_n_32_12),.A2(multiplier_0_n_32_28),.ZN(multiplier_0_n_32_398));
	OR3_X1_LVT multiplier_0i_32_372 (.A1(multiplier_0_n_32_396),.A2(multiplier_0_n_32_397),.A3(multiplier_0_n_32_398),.ZN(multiplier_0_n_32_395));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b8___05F05d (.D(multiplier_0_per_din_msk[8]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[8]),.QN());
	NAND2_X1_LVT multiplier_0i_32_76 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_32_76));
	NAND2_X1_LVT multiplier_0i_32_92 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_32_92));
	NOR2_X1_LVT multiplier_0i_32_366 (.A1(multiplier_0_n_32_76),.A2(multiplier_0_n_32_92),.ZN(multiplier_0_n_32_389));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b9___05F05d (.D(multiplier_0_per_din_msk[9]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[9]),.QN());
	NAND2_X1_LVT multiplier_0i_32_60 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_32_60));
	NOR2_X1_LVT multiplier_0i_32_367 (.A1(multiplier_0_n_32_60),.A2(multiplier_0_n_32_92),.ZN(multiplier_0_n_32_390));
	NOR2_X1_LVT multiplier_0i_32_368 (.A1(multiplier_0_n_32_60),.A2(multiplier_0_n_32_76),.ZN(multiplier_0_n_32_391));
	OR3_X1_LVT multiplier_0i_32_365 (.A1(multiplier_0_n_32_389),.A2(multiplier_0_n_32_390),.A3(multiplier_0_n_32_391),.ZN(multiplier_0_n_32_388));
	NAND2_X1_LVT multiplier_0i_32_140 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_32_140));
	NAND2_X1_LVT multiplier_0i_32_124 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_32_124));
	INV_X1_LVT multiplier_0i_32_358 (.A(multiplier_0_n_32_124),.ZN(multiplier_0_n_32_381));
	NAND2_X1_LVT multiplier_0i_32_357 (.A1(multiplier_0_n_32_140),.A2(multiplier_0_n_32_381),.ZN(multiplier_0_n_32_380));
	NAND2_X1_LVT multiplier_0i_32_108 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_32_108));
	INV_X1_LVT multiplier_0i_32_360 (.A(multiplier_0_n_32_108),.ZN(multiplier_0_n_32_383));
	NAND2_X1_LVT multiplier_0i_32_359 (.A1(multiplier_0_n_32_140),.A2(multiplier_0_n_32_383),.ZN(multiplier_0_n_32_382));
	OR2_X1_LVT multiplier_0i_32_361 (.A1(multiplier_0_n_32_108),.A2(multiplier_0_n_32_124),.ZN(multiplier_0_n_32_384));
	NAND3_X1_LVT multiplier_0i_32_356 (.A1(multiplier_0_n_32_380),.A2(multiplier_0_n_32_382),.A3(multiplier_0_n_32_384),.ZN(multiplier_0_n_32_379));
	FA_X1_LVT multiplier_0i_32_402 (.A(multiplier_0_n_32_395),.B(multiplier_0_n_32_388),.CI(multiplier_0_n_32_379),.CO(multiplier_0_n_32_430),.S(multiplier_0_n_32_429));
	NAND2_X1_LVT multiplier_0i_32_26 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_32_26));
	NAND2_X1_LVT multiplier_0i_32_42 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_32_42));
	NOR2_X1_LVT multiplier_0i_32_321 (.A1(multiplier_0_n_32_26),.A2(multiplier_0_n_32_42),.ZN(multiplier_0_n_32_336));
	NAND2_X1_LVT multiplier_0i_32_10 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_32_10));
	NOR2_X1_LVT multiplier_0i_32_322 (.A1(multiplier_0_n_32_10),.A2(multiplier_0_n_32_42),.ZN(multiplier_0_n_32_337));
	NOR2_X1_LVT multiplier_0i_32_323 (.A1(multiplier_0_n_32_10),.A2(multiplier_0_n_32_26),.ZN(multiplier_0_n_32_338));
	OR3_X1_LVT multiplier_0i_32_320 (.A1(multiplier_0_n_32_336),.A2(multiplier_0_n_32_337),.A3(multiplier_0_n_32_338),.ZN(multiplier_0_n_32_335));
	NAND2_X1_LVT multiplier_0i_32_74 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_32_74));
	NAND2_X1_LVT multiplier_0i_32_90 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_32_90));
	NOR2_X1_LVT multiplier_0i_32_314 (.A1(multiplier_0_n_32_74),.A2(multiplier_0_n_32_90),.ZN(multiplier_0_n_32_329));
	NAND2_X1_LVT multiplier_0i_32_58 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_32_58));
	NOR2_X1_LVT multiplier_0i_32_315 (.A1(multiplier_0_n_32_58),.A2(multiplier_0_n_32_90),.ZN(multiplier_0_n_32_330));
	NOR2_X1_LVT multiplier_0i_32_316 (.A1(multiplier_0_n_32_58),.A2(multiplier_0_n_32_74),.ZN(multiplier_0_n_32_331));
	OR3_X1_LVT multiplier_0i_32_313 (.A1(multiplier_0_n_32_329),.A2(multiplier_0_n_32_330),.A3(multiplier_0_n_32_331),.ZN(multiplier_0_n_32_328));
	NAND2_X1_LVT multiplier_0i_32_138 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_32_138));
	NAND2_X1_LVT multiplier_0i_32_122 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_32_122));
	INV_X1_LVT multiplier_0i_32_306 (.A(multiplier_0_n_32_122),.ZN(multiplier_0_n_32_321));
	NAND2_X1_LVT multiplier_0i_32_305 (.A1(multiplier_0_n_32_138),.A2(multiplier_0_n_32_321),.ZN(multiplier_0_n_32_320));
	NAND2_X1_LVT multiplier_0i_32_106 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_32_106));
	INV_X1_LVT multiplier_0i_32_308 (.A(multiplier_0_n_32_106),.ZN(multiplier_0_n_32_323));
	NAND2_X1_LVT multiplier_0i_32_307 (.A1(multiplier_0_n_32_138),.A2(multiplier_0_n_32_323),.ZN(multiplier_0_n_32_322));
	OR2_X1_LVT multiplier_0i_32_309 (.A1(multiplier_0_n_32_106),.A2(multiplier_0_n_32_122),.ZN(multiplier_0_n_32_324));
	NAND3_X1_LVT multiplier_0i_32_304 (.A1(multiplier_0_n_32_320),.A2(multiplier_0_n_32_322),.A3(multiplier_0_n_32_324),.ZN(multiplier_0_n_32_319));
	FA_X1_LVT multiplier_0i_32_350 (.A(multiplier_0_n_32_335),.B(multiplier_0_n_32_328),.CI(multiplier_0_n_32_319),.CO(multiplier_0_n_32_370),.S(multiplier_0_n_32_369));
	XNOR2_X1_LVT multiplier_0i_32_369 (.A(multiplier_0_n_32_44),.B(multiplier_0_n_32_28),.ZN(multiplier_0_n_32_392));
	XNOR2_X1_LVT multiplier_0i_32_370 (.A(multiplier_0_n_32_392),.B(multiplier_0_n_32_12),.ZN(multiplier_0_n_32_393));
	INV_X1_LVT multiplier_0i_32_371 (.A(multiplier_0_n_32_393),.ZN(multiplier_0_n_32_394));
	XNOR2_X1_LVT multiplier_0i_32_362 (.A(multiplier_0_n_32_92),.B(multiplier_0_n_32_76),.ZN(multiplier_0_n_32_385));
	XNOR2_X1_LVT multiplier_0i_32_363 (.A(multiplier_0_n_32_385),.B(multiplier_0_n_32_60),.ZN(multiplier_0_n_32_386));
	INV_X1_LVT multiplier_0i_32_364 (.A(multiplier_0_n_32_386),.ZN(multiplier_0_n_32_387));
	FA_X1_LVT multiplier_0i_32_377 (.A(multiplier_0_n_32_370),.B(multiplier_0_n_32_394),.CI(multiplier_0_n_32_387),.CO(multiplier_0_n_32_402),.S(multiplier_0_n_32_401));
	FA_X1_LVT multiplier_0i_32_404 (.A(multiplier_0_n_32_408),.B(multiplier_0_n_32_429),.CI(multiplier_0_n_32_402),.CO(multiplier_0_n_32_434),.S(multiplier_0_n_32_433));
	NAND2_X1_LVT multiplier_0i_32_46 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_32_46));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b13___05F05d (.D(multiplier_0_per_din_msk[13]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[13]),.QN());
	NAND2_X1_LVT multiplier_0i_32_30 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_32_30));
	XNOR2_X1_LVT multiplier_0i_32_421 (.A(multiplier_0_n_32_46),.B(multiplier_0_n_32_30),.ZN(multiplier_0_n_32_452));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b14___05F05d (.D(multiplier_0_per_din_msk[14]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[14]),.QN());
	NAND2_X1_LVT multiplier_0i_32_14 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_32_14));
	XNOR2_X1_LVT multiplier_0i_32_422 (.A(multiplier_0_n_32_452),.B(multiplier_0_n_32_14),.ZN(multiplier_0_n_32_453));
	INV_X1_LVT multiplier_0i_32_423 (.A(multiplier_0_n_32_453),.ZN(multiplier_0_n_32_454));
	NAND2_X1_LVT multiplier_0i_32_94 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_32_94));
	NAND2_X1_LVT multiplier_0i_32_78 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_32_78));
	XNOR2_X1_LVT multiplier_0i_32_414 (.A(multiplier_0_n_32_94),.B(multiplier_0_n_32_78),.ZN(multiplier_0_n_32_445));
	NAND2_X1_LVT multiplier_0i_32_62 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_32_62));
	XNOR2_X1_LVT multiplier_0i_32_415 (.A(multiplier_0_n_32_445),.B(multiplier_0_n_32_62),.ZN(multiplier_0_n_32_446));
	INV_X1_LVT multiplier_0i_32_416 (.A(multiplier_0_n_32_446),.ZN(multiplier_0_n_32_447));
	FA_X1_LVT multiplier_0i_32_429 (.A(multiplier_0_n_32_430),.B(multiplier_0_n_32_454),.CI(multiplier_0_n_32_447),.CO(multiplier_0_n_32_462),.S(multiplier_0_n_32_461));
	NAND2_X1_LVT multiplier_0i_32_142 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_32_142));
	NAND2_X1_LVT multiplier_0i_32_126 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_32_126));
	XNOR2_X1_LVT multiplier_0i_32_406 (.A(multiplier_0_n_32_142),.B(multiplier_0_n_32_126),.ZN(multiplier_0_n_32_437));
	NAND2_X1_LVT multiplier_0i_32_110 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_32_110));
	XNOR2_X1_LVT multiplier_0i_32_407 (.A(multiplier_0_n_32_437),.B(multiplier_0_n_32_110),.ZN(multiplier_0_n_32_438));
	NAND2_X1_LVT multiplier_0i_32_29 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_32_29));
	NAND2_X1_LVT multiplier_0i_32_45 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_32_45));
	NOR2_X1_LVT multiplier_0i_32_399 (.A1(multiplier_0_n_32_29),.A2(multiplier_0_n_32_45),.ZN(multiplier_0_n_32_426));
	NAND2_X1_LVT multiplier_0i_32_13 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_32_13));
	NOR2_X1_LVT multiplier_0i_32_400 (.A1(multiplier_0_n_32_13),.A2(multiplier_0_n_32_45),.ZN(multiplier_0_n_32_427));
	NOR2_X1_LVT multiplier_0i_32_401 (.A1(multiplier_0_n_32_13),.A2(multiplier_0_n_32_29),.ZN(multiplier_0_n_32_428));
	OR3_X1_LVT multiplier_0i_32_398 (.A1(multiplier_0_n_32_426),.A2(multiplier_0_n_32_427),.A3(multiplier_0_n_32_428),.ZN(multiplier_0_n_32_425));
	NAND2_X1_LVT multiplier_0i_32_77 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_32_77));
	NAND2_X1_LVT multiplier_0i_32_93 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_32_93));
	NOR2_X1_LVT multiplier_0i_32_392 (.A1(multiplier_0_n_32_77),.A2(multiplier_0_n_32_93),.ZN(multiplier_0_n_32_419));
	NAND2_X1_LVT multiplier_0i_32_61 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_32_61));
	NOR2_X1_LVT multiplier_0i_32_393 (.A1(multiplier_0_n_32_61),.A2(multiplier_0_n_32_93),.ZN(multiplier_0_n_32_420));
	NOR2_X1_LVT multiplier_0i_32_394 (.A1(multiplier_0_n_32_61),.A2(multiplier_0_n_32_77),.ZN(multiplier_0_n_32_421));
	OR3_X1_LVT multiplier_0i_32_391 (.A1(multiplier_0_n_32_419),.A2(multiplier_0_n_32_420),.A3(multiplier_0_n_32_421),.ZN(multiplier_0_n_32_418));
	INV_X1_LVT multiplier_0i_32_384 (.A(multiplier_0_n_32_125),.ZN(multiplier_0_n_32_411));
	NAND2_X1_LVT multiplier_0i_32_383 (.A1(multiplier_0_n_32_141),.A2(multiplier_0_n_32_411),.ZN(multiplier_0_n_32_410));
	INV_X1_LVT multiplier_0i_32_386 (.A(multiplier_0_n_32_109),.ZN(multiplier_0_n_32_413));
	NAND2_X1_LVT multiplier_0i_32_385 (.A1(multiplier_0_n_32_141),.A2(multiplier_0_n_32_413),.ZN(multiplier_0_n_32_412));
	OR2_X1_LVT multiplier_0i_32_387 (.A1(multiplier_0_n_32_109),.A2(multiplier_0_n_32_125),.ZN(multiplier_0_n_32_414));
	NAND3_X1_LVT multiplier_0i_32_382 (.A1(multiplier_0_n_32_410),.A2(multiplier_0_n_32_412),.A3(multiplier_0_n_32_414),.ZN(multiplier_0_n_32_409));
	FA_X1_LVT multiplier_0i_32_428 (.A(multiplier_0_n_32_425),.B(multiplier_0_n_32_418),.CI(multiplier_0_n_32_409),.CO(multiplier_0_n_32_460),.S(multiplier_0_n_32_459));
	NAND2_X1_LVT multiplier_0i_32_27 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_32_27));
	NAND2_X1_LVT multiplier_0i_32_43 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_32_43));
	NOR2_X1_LVT multiplier_0i_32_347 (.A1(multiplier_0_n_32_27),.A2(multiplier_0_n_32_43),.ZN(multiplier_0_n_32_366));
	NAND2_X1_LVT multiplier_0i_32_11 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_32_11));
	NOR2_X1_LVT multiplier_0i_32_348 (.A1(multiplier_0_n_32_11),.A2(multiplier_0_n_32_43),.ZN(multiplier_0_n_32_367));
	NOR2_X1_LVT multiplier_0i_32_349 (.A1(multiplier_0_n_32_11),.A2(multiplier_0_n_32_27),.ZN(multiplier_0_n_32_368));
	OR3_X1_LVT multiplier_0i_32_346 (.A1(multiplier_0_n_32_366),.A2(multiplier_0_n_32_367),.A3(multiplier_0_n_32_368),.ZN(multiplier_0_n_32_365));
	NAND2_X1_LVT multiplier_0i_32_75 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_32_75));
	NAND2_X1_LVT multiplier_0i_32_91 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_32_91));
	NOR2_X1_LVT multiplier_0i_32_340 (.A1(multiplier_0_n_32_75),.A2(multiplier_0_n_32_91),.ZN(multiplier_0_n_32_359));
	NAND2_X1_LVT multiplier_0i_32_59 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_32_59));
	NOR2_X1_LVT multiplier_0i_32_341 (.A1(multiplier_0_n_32_59),.A2(multiplier_0_n_32_91),.ZN(multiplier_0_n_32_360));
	NOR2_X1_LVT multiplier_0i_32_342 (.A1(multiplier_0_n_32_59),.A2(multiplier_0_n_32_75),.ZN(multiplier_0_n_32_361));
	OR3_X1_LVT multiplier_0i_32_339 (.A1(multiplier_0_n_32_359),.A2(multiplier_0_n_32_360),.A3(multiplier_0_n_32_361),.ZN(multiplier_0_n_32_358));
	NAND2_X1_LVT multiplier_0i_32_139 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_32_139));
	NAND2_X1_LVT multiplier_0i_32_123 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_32_123));
	INV_X1_LVT multiplier_0i_32_332 (.A(multiplier_0_n_32_123),.ZN(multiplier_0_n_32_351));
	NAND2_X1_LVT multiplier_0i_32_331 (.A1(multiplier_0_n_32_139),.A2(multiplier_0_n_32_351),.ZN(multiplier_0_n_32_350));
	NAND2_X1_LVT multiplier_0i_32_107 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_32_107));
	INV_X1_LVT multiplier_0i_32_334 (.A(multiplier_0_n_32_107),.ZN(multiplier_0_n_32_353));
	NAND2_X1_LVT multiplier_0i_32_333 (.A1(multiplier_0_n_32_139),.A2(multiplier_0_n_32_353),.ZN(multiplier_0_n_32_352));
	OR2_X1_LVT multiplier_0i_32_335 (.A1(multiplier_0_n_32_107),.A2(multiplier_0_n_32_123),.ZN(multiplier_0_n_32_354));
	NAND3_X1_LVT multiplier_0i_32_330 (.A1(multiplier_0_n_32_350),.A2(multiplier_0_n_32_352),.A3(multiplier_0_n_32_354),.ZN(multiplier_0_n_32_349));
	FA_X1_LVT multiplier_0i_32_376 (.A(multiplier_0_n_32_365),.B(multiplier_0_n_32_358),.CI(multiplier_0_n_32_349),.CO(multiplier_0_n_32_400),.S(multiplier_0_n_32_399));
	XNOR2_X1_LVT multiplier_0i_32_395 (.A(multiplier_0_n_32_45),.B(multiplier_0_n_32_29),.ZN(multiplier_0_n_32_422));
	XNOR2_X1_LVT multiplier_0i_32_396 (.A(multiplier_0_n_32_422),.B(multiplier_0_n_32_13),.ZN(multiplier_0_n_32_423));
	INV_X1_LVT multiplier_0i_32_397 (.A(multiplier_0_n_32_423),.ZN(multiplier_0_n_32_424));
	XNOR2_X1_LVT multiplier_0i_32_388 (.A(multiplier_0_n_32_93),.B(multiplier_0_n_32_77),.ZN(multiplier_0_n_32_415));
	XNOR2_X1_LVT multiplier_0i_32_389 (.A(multiplier_0_n_32_415),.B(multiplier_0_n_32_61),.ZN(multiplier_0_n_32_416));
	INV_X1_LVT multiplier_0i_32_390 (.A(multiplier_0_n_32_416),.ZN(multiplier_0_n_32_417));
	FA_X1_LVT multiplier_0i_32_403 (.A(multiplier_0_n_32_400),.B(multiplier_0_n_32_424),.CI(multiplier_0_n_32_417),.CO(multiplier_0_n_32_432),.S(multiplier_0_n_32_431));
	FA_X1_LVT multiplier_0i_32_430 (.A(multiplier_0_n_32_438),.B(multiplier_0_n_32_459),.CI(multiplier_0_n_32_432),.CO(multiplier_0_n_32_464),.S(multiplier_0_n_32_463));
	FA_X1_LVT multiplier_0i_32_431 (.A(multiplier_0_n_32_434),.B(multiplier_0_n_32_461),.CI(multiplier_0_n_32_463),.CO(multiplier_0_n_32_466),.S(multiplier_0_n_32_465));
	NAND2_X1_LVT multiplier_0i_32_47 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_32_47));
	NAND2_X1_LVT multiplier_0i_32_31 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_32_31));
	XNOR2_X1_LVT multiplier_0i_32_447 (.A(multiplier_0_n_32_47),.B(multiplier_0_n_32_31),.ZN(multiplier_0_n_32_482));
	DFFR_X1_LVT multiplier_0op1_reg___05F05b15___05F05d (.D(multiplier_0_per_din_msk[15]),.RN(multiplier_0_n_38),.CK(multiplier_0_n_41),.Q(multiplier_0_op1[15]),.QN());
	NAND2_X1_LVT multiplier_0i_32_15 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_32_15));
	XNOR2_X1_LVT multiplier_0i_32_448 (.A(multiplier_0_n_32_482),.B(multiplier_0_n_32_15),.ZN(multiplier_0_n_32_483));
	INV_X1_LVT multiplier_0i_32_449 (.A(multiplier_0_n_32_483),.ZN(multiplier_0_n_32_484));
	NAND2_X1_LVT multiplier_0i_32_95 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_32_95));
	NAND2_X1_LVT multiplier_0i_32_79 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_32_79));
	XNOR2_X1_LVT multiplier_0i_32_440 (.A(multiplier_0_n_32_95),.B(multiplier_0_n_32_79),.ZN(multiplier_0_n_32_475));
	NAND2_X1_LVT multiplier_0i_32_63 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_32_63));
	XNOR2_X1_LVT multiplier_0i_32_441 (.A(multiplier_0_n_32_475),.B(multiplier_0_n_32_63),.ZN(multiplier_0_n_32_476));
	INV_X1_LVT multiplier_0i_32_442 (.A(multiplier_0_n_32_476),.ZN(multiplier_0_n_32_477));
	FA_X1_LVT multiplier_0i_32_455 (.A(multiplier_0_n_32_460),.B(multiplier_0_n_32_484),.CI(multiplier_0_n_32_477),.CO(multiplier_0_n_32_492),.S(multiplier_0_n_32_491));
	NAND2_X1_LVT multiplier_0i_32_143 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_32_143));
	NAND2_X1_LVT multiplier_0i_32_127 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_32_127));
	XNOR2_X1_LVT multiplier_0i_32_432 (.A(multiplier_0_n_32_143),.B(multiplier_0_n_32_127),.ZN(multiplier_0_n_32_467));
	NAND2_X1_LVT multiplier_0i_32_111 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_32_111));
	XNOR2_X1_LVT multiplier_0i_32_433 (.A(multiplier_0_n_32_467),.B(multiplier_0_n_32_111),.ZN(multiplier_0_n_32_468));
	NOR2_X1_LVT multiplier_0i_32_425 (.A1(multiplier_0_n_32_30),.A2(multiplier_0_n_32_46),.ZN(multiplier_0_n_32_456));
	NOR2_X1_LVT multiplier_0i_32_426 (.A1(multiplier_0_n_32_14),.A2(multiplier_0_n_32_46),.ZN(multiplier_0_n_32_457));
	NOR2_X1_LVT multiplier_0i_32_427 (.A1(multiplier_0_n_32_14),.A2(multiplier_0_n_32_30),.ZN(multiplier_0_n_32_458));
	OR3_X1_LVT multiplier_0i_32_424 (.A1(multiplier_0_n_32_456),.A2(multiplier_0_n_32_457),.A3(multiplier_0_n_32_458),.ZN(multiplier_0_n_32_455));
	NOR2_X1_LVT multiplier_0i_32_418 (.A1(multiplier_0_n_32_78),.A2(multiplier_0_n_32_94),.ZN(multiplier_0_n_32_449));
	NOR2_X1_LVT multiplier_0i_32_419 (.A1(multiplier_0_n_32_62),.A2(multiplier_0_n_32_94),.ZN(multiplier_0_n_32_450));
	NOR2_X1_LVT multiplier_0i_32_420 (.A1(multiplier_0_n_32_62),.A2(multiplier_0_n_32_78),.ZN(multiplier_0_n_32_451));
	OR3_X1_LVT multiplier_0i_32_417 (.A1(multiplier_0_n_32_449),.A2(multiplier_0_n_32_450),.A3(multiplier_0_n_32_451),.ZN(multiplier_0_n_32_448));
	INV_X1_LVT multiplier_0i_32_410 (.A(multiplier_0_n_32_126),.ZN(multiplier_0_n_32_441));
	NAND2_X1_LVT multiplier_0i_32_409 (.A1(multiplier_0_n_32_142),.A2(multiplier_0_n_32_441),.ZN(multiplier_0_n_32_440));
	INV_X1_LVT multiplier_0i_32_412 (.A(multiplier_0_n_32_110),.ZN(multiplier_0_n_32_443));
	NAND2_X1_LVT multiplier_0i_32_411 (.A1(multiplier_0_n_32_142),.A2(multiplier_0_n_32_443),.ZN(multiplier_0_n_32_442));
	OR2_X1_LVT multiplier_0i_32_413 (.A1(multiplier_0_n_32_110),.A2(multiplier_0_n_32_126),.ZN(multiplier_0_n_32_444));
	NAND3_X1_LVT multiplier_0i_32_408 (.A1(multiplier_0_n_32_440),.A2(multiplier_0_n_32_442),.A3(multiplier_0_n_32_444),.ZN(multiplier_0_n_32_439));
	FA_X1_LVT multiplier_0i_32_454 (.A(multiplier_0_n_32_455),.B(multiplier_0_n_32_448),.CI(multiplier_0_n_32_439),.CO(multiplier_0_n_32_490),.S(multiplier_0_n_32_489));
	FA_X1_LVT multiplier_0i_32_456 (.A(multiplier_0_n_32_468),.B(multiplier_0_n_32_489),.CI(multiplier_0_n_32_462),.CO(multiplier_0_n_32_494),.S(multiplier_0_n_32_493));
	FA_X1_LVT multiplier_0i_32_457 (.A(multiplier_0_n_32_464),.B(multiplier_0_n_32_491),.CI(multiplier_0_n_32_493),.CO(multiplier_0_n_32_496),.S(multiplier_0_n_32_495));
	XNOR2_X1_LVT multiplier_0i_32_354 (.A(multiplier_0_n_32_140),.B(multiplier_0_n_32_124),.ZN(multiplier_0_n_32_377));
	XNOR2_X1_LVT multiplier_0i_32_355 (.A(multiplier_0_n_32_377),.B(multiplier_0_n_32_108),.ZN(multiplier_0_n_32_378));
	NAND2_X1_LVT multiplier_0i_32_25 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_32_25));
	NAND2_X1_LVT multiplier_0i_32_41 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_32_41));
	NOR2_X1_LVT multiplier_0i_32_295 (.A1(multiplier_0_n_32_25),.A2(multiplier_0_n_32_41),.ZN(multiplier_0_n_32_306));
	NAND2_X1_LVT multiplier_0i_32_9 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_32_9));
	NOR2_X1_LVT multiplier_0i_32_296 (.A1(multiplier_0_n_32_9),.A2(multiplier_0_n_32_41),.ZN(multiplier_0_n_32_307));
	NOR2_X1_LVT multiplier_0i_32_297 (.A1(multiplier_0_n_32_9),.A2(multiplier_0_n_32_25),.ZN(multiplier_0_n_32_308));
	OR3_X1_LVT multiplier_0i_32_294 (.A1(multiplier_0_n_32_306),.A2(multiplier_0_n_32_307),.A3(multiplier_0_n_32_308),.ZN(multiplier_0_n_32_305));
	NAND2_X1_LVT multiplier_0i_32_73 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_32_73));
	NAND2_X1_LVT multiplier_0i_32_89 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_32_89));
	NOR2_X1_LVT multiplier_0i_32_288 (.A1(multiplier_0_n_32_73),.A2(multiplier_0_n_32_89),.ZN(multiplier_0_n_32_299));
	NAND2_X1_LVT multiplier_0i_32_57 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_32_57));
	NOR2_X1_LVT multiplier_0i_32_289 (.A1(multiplier_0_n_32_57),.A2(multiplier_0_n_32_89),.ZN(multiplier_0_n_32_300));
	NOR2_X1_LVT multiplier_0i_32_290 (.A1(multiplier_0_n_32_57),.A2(multiplier_0_n_32_73),.ZN(multiplier_0_n_32_301));
	OR3_X1_LVT multiplier_0i_32_287 (.A1(multiplier_0_n_32_299),.A2(multiplier_0_n_32_300),.A3(multiplier_0_n_32_301),.ZN(multiplier_0_n_32_298));
	NAND2_X1_LVT multiplier_0i_32_137 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_32_137));
	NAND2_X1_LVT multiplier_0i_32_121 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_32_121));
	INV_X1_LVT multiplier_0i_32_280 (.A(multiplier_0_n_32_121),.ZN(multiplier_0_n_32_291));
	NAND2_X1_LVT multiplier_0i_32_279 (.A1(multiplier_0_n_32_137),.A2(multiplier_0_n_32_291),.ZN(multiplier_0_n_32_290));
	NAND2_X1_LVT multiplier_0i_32_105 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_32_105));
	INV_X1_LVT multiplier_0i_32_282 (.A(multiplier_0_n_32_105),.ZN(multiplier_0_n_32_293));
	NAND2_X1_LVT multiplier_0i_32_281 (.A1(multiplier_0_n_32_137),.A2(multiplier_0_n_32_293),.ZN(multiplier_0_n_32_292));
	OR2_X1_LVT multiplier_0i_32_283 (.A1(multiplier_0_n_32_105),.A2(multiplier_0_n_32_121),.ZN(multiplier_0_n_32_294));
	NAND3_X1_LVT multiplier_0i_32_278 (.A1(multiplier_0_n_32_290),.A2(multiplier_0_n_32_292),.A3(multiplier_0_n_32_294),.ZN(multiplier_0_n_32_289));
	FA_X1_LVT multiplier_0i_32_324 (.A(multiplier_0_n_32_305),.B(multiplier_0_n_32_298),.CI(multiplier_0_n_32_289),.CO(multiplier_0_n_32_340),.S(multiplier_0_n_32_339));
	XNOR2_X1_LVT multiplier_0i_32_343 (.A(multiplier_0_n_32_43),.B(multiplier_0_n_32_27),.ZN(multiplier_0_n_32_362));
	XNOR2_X1_LVT multiplier_0i_32_344 (.A(multiplier_0_n_32_362),.B(multiplier_0_n_32_11),.ZN(multiplier_0_n_32_363));
	INV_X1_LVT multiplier_0i_32_345 (.A(multiplier_0_n_32_363),.ZN(multiplier_0_n_32_364));
	XNOR2_X1_LVT multiplier_0i_32_336 (.A(multiplier_0_n_32_91),.B(multiplier_0_n_32_75),.ZN(multiplier_0_n_32_355));
	XNOR2_X1_LVT multiplier_0i_32_337 (.A(multiplier_0_n_32_355),.B(multiplier_0_n_32_59),.ZN(multiplier_0_n_32_356));
	INV_X1_LVT multiplier_0i_32_338 (.A(multiplier_0_n_32_356),.ZN(multiplier_0_n_32_357));
	FA_X1_LVT multiplier_0i_32_351 (.A(multiplier_0_n_32_340),.B(multiplier_0_n_32_364),.CI(multiplier_0_n_32_357),.CO(multiplier_0_n_32_372),.S(multiplier_0_n_32_371));
	FA_X1_LVT multiplier_0i_32_378 (.A(multiplier_0_n_32_378),.B(multiplier_0_n_32_399),.CI(multiplier_0_n_32_372),.CO(multiplier_0_n_32_404),.S(multiplier_0_n_32_403));
	FA_X1_LVT multiplier_0i_32_405 (.A(multiplier_0_n_32_404),.B(multiplier_0_n_32_431),.CI(multiplier_0_n_32_433),.CO(multiplier_0_n_32_436),.S(multiplier_0_n_32_435));
	XNOR2_X1_LVT multiplier_0i_32_328 (.A(multiplier_0_n_32_139),.B(multiplier_0_n_32_123),.ZN(multiplier_0_n_32_347));
	XNOR2_X1_LVT multiplier_0i_32_329 (.A(multiplier_0_n_32_347),.B(multiplier_0_n_32_107),.ZN(multiplier_0_n_32_348));
	NAND2_X1_LVT multiplier_0i_32_40 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_32_40));
	NAND2_X1_LVT multiplier_0i_32_56 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_32_56));
	NOR2_X1_LVT multiplier_0i_32_262 (.A1(multiplier_0_n_32_40),.A2(multiplier_0_n_32_56),.ZN(multiplier_0_n_32_270));
	NAND2_X1_LVT multiplier_0i_32_24 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_32_24));
	NOR2_X1_LVT multiplier_0i_32_263 (.A1(multiplier_0_n_32_24),.A2(multiplier_0_n_32_56),.ZN(multiplier_0_n_32_271));
	NOR2_X1_LVT multiplier_0i_32_264 (.A1(multiplier_0_n_32_24),.A2(multiplier_0_n_32_40),.ZN(multiplier_0_n_32_272));
	OR3_X1_LVT multiplier_0i_32_261 (.A1(multiplier_0_n_32_270),.A2(multiplier_0_n_32_271),.A3(multiplier_0_n_32_272),.ZN(multiplier_0_n_32_269));
	NAND2_X1_LVT multiplier_0i_32_88 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_32_88));
	NAND2_X1_LVT multiplier_0i_32_104 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_32_104));
	NOR2_X1_LVT multiplier_0i_32_255 (.A1(multiplier_0_n_32_88),.A2(multiplier_0_n_32_104),.ZN(multiplier_0_n_32_263));
	NAND2_X1_LVT multiplier_0i_32_72 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_32_72));
	NOR2_X1_LVT multiplier_0i_32_256 (.A1(multiplier_0_n_32_72),.A2(multiplier_0_n_32_104),.ZN(multiplier_0_n_32_264));
	NOR2_X1_LVT multiplier_0i_32_257 (.A1(multiplier_0_n_32_72),.A2(multiplier_0_n_32_88),.ZN(multiplier_0_n_32_265));
	OR3_X1_LVT multiplier_0i_32_254 (.A1(multiplier_0_n_32_263),.A2(multiplier_0_n_32_264),.A3(multiplier_0_n_32_265),.ZN(multiplier_0_n_32_262));
	NAND2_X1_LVT multiplier_0i_32_120 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_32_120));
	NAND2_X1_LVT multiplier_0i_32_136 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[0]),.ZN(multiplier_0_n_32_136));
	INV_X1_LVT multiplier_0i_32_250 (.A(multiplier_0_n_32_136),.ZN(multiplier_0_n_32_258));
	NAND2_X1_LVT multiplier_0i_32_249 (.A1(multiplier_0_n_32_120),.A2(multiplier_0_n_32_258),.ZN(multiplier_0_n_32_257));
	FA_X1_LVT multiplier_0i_32_298 (.A(multiplier_0_n_32_269),.B(multiplier_0_n_32_262),.CI(multiplier_0_n_32_257),.CO(multiplier_0_n_32_310),.S(multiplier_0_n_32_309));
	XNOR2_X1_LVT multiplier_0i_32_317 (.A(multiplier_0_n_32_42),.B(multiplier_0_n_32_26),.ZN(multiplier_0_n_32_332));
	XNOR2_X1_LVT multiplier_0i_32_318 (.A(multiplier_0_n_32_332),.B(multiplier_0_n_32_10),.ZN(multiplier_0_n_32_333));
	INV_X1_LVT multiplier_0i_32_319 (.A(multiplier_0_n_32_333),.ZN(multiplier_0_n_32_334));
	XNOR2_X1_LVT multiplier_0i_32_310 (.A(multiplier_0_n_32_90),.B(multiplier_0_n_32_74),.ZN(multiplier_0_n_32_325));
	XNOR2_X1_LVT multiplier_0i_32_311 (.A(multiplier_0_n_32_325),.B(multiplier_0_n_32_58),.ZN(multiplier_0_n_32_326));
	INV_X1_LVT multiplier_0i_32_312 (.A(multiplier_0_n_32_326),.ZN(multiplier_0_n_32_327));
	FA_X1_LVT multiplier_0i_32_325 (.A(multiplier_0_n_32_310),.B(multiplier_0_n_32_334),.CI(multiplier_0_n_32_327),.CO(multiplier_0_n_32_342),.S(multiplier_0_n_32_341));
	FA_X1_LVT multiplier_0i_32_352 (.A(multiplier_0_n_32_348),.B(multiplier_0_n_32_369),.CI(multiplier_0_n_32_342),.CO(multiplier_0_n_32_374),.S(multiplier_0_n_32_373));
	FA_X1_LVT multiplier_0i_32_379 (.A(multiplier_0_n_32_374),.B(multiplier_0_n_32_401),.CI(multiplier_0_n_32_403),.CO(multiplier_0_n_32_406),.S(multiplier_0_n_32_405));
	XNOR2_X1_LVT multiplier_0i_32_302 (.A(multiplier_0_n_32_138),.B(multiplier_0_n_32_122),.ZN(multiplier_0_n_32_317));
	XNOR2_X1_LVT multiplier_0i_32_303 (.A(multiplier_0_n_32_317),.B(multiplier_0_n_32_106),.ZN(multiplier_0_n_32_318));
	NOR2_X1_LVT multiplier_0i_32_233 (.A1(multiplier_0_n_32_55),.A2(multiplier_0_n_32_71),.ZN(multiplier_0_n_32_238));
	NOR2_X1_LVT multiplier_0i_32_234 (.A1(multiplier_0_n_32_39),.A2(multiplier_0_n_32_71),.ZN(multiplier_0_n_32_239));
	NOR2_X1_LVT multiplier_0i_32_235 (.A1(multiplier_0_n_32_39),.A2(multiplier_0_n_32_55),.ZN(multiplier_0_n_32_240));
	OR3_X1_LVT multiplier_0i_32_232 (.A1(multiplier_0_n_32_238),.A2(multiplier_0_n_32_239),.A3(multiplier_0_n_32_240),.ZN(multiplier_0_n_32_237));
	NAND2_X1_LVT multiplier_0i_32_8 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_32_8));
	INV_X1_LVT multiplier_0i_32_270 (.A(multiplier_0_n_32_8),.ZN(multiplier_0_n_32_278));
	NAND2_X1_LVT multiplier_0i_32_269 (.A1(multiplier_0_n_32_237),.A2(multiplier_0_n_32_278),.ZN(multiplier_0_n_32_277));
	NOR2_X1_LVT multiplier_0i_32_226 (.A1(multiplier_0_n_32_103),.A2(multiplier_0_n_32_119),.ZN(multiplier_0_n_32_231));
	NOR2_X1_LVT multiplier_0i_32_227 (.A1(multiplier_0_n_32_87),.A2(multiplier_0_n_32_119),.ZN(multiplier_0_n_32_232));
	NOR2_X1_LVT multiplier_0i_32_228 (.A1(multiplier_0_n_32_87),.A2(multiplier_0_n_32_103),.ZN(multiplier_0_n_32_233));
	OR3_X1_LVT multiplier_0i_32_225 (.A1(multiplier_0_n_32_231),.A2(multiplier_0_n_32_232),.A3(multiplier_0_n_32_233),.ZN(multiplier_0_n_32_230));
	NAND2_X1_LVT multiplier_0i_32_271 (.A1(multiplier_0_n_32_230),.A2(multiplier_0_n_32_278),.ZN(multiplier_0_n_32_279));
	NAND2_X1_LVT multiplier_0i_32_272 (.A1(multiplier_0_n_32_230),.A2(multiplier_0_n_32_237),.ZN(multiplier_0_n_32_280));
	NAND3_X1_LVT multiplier_0i_32_268 (.A1(multiplier_0_n_32_277),.A2(multiplier_0_n_32_279),.A3(multiplier_0_n_32_280),.ZN(multiplier_0_n_32_276));
	XNOR2_X1_LVT multiplier_0i_32_291 (.A(multiplier_0_n_32_41),.B(multiplier_0_n_32_25),.ZN(multiplier_0_n_32_302));
	XNOR2_X1_LVT multiplier_0i_32_292 (.A(multiplier_0_n_32_302),.B(multiplier_0_n_32_9),.ZN(multiplier_0_n_32_303));
	INV_X1_LVT multiplier_0i_32_293 (.A(multiplier_0_n_32_303),.ZN(multiplier_0_n_32_304));
	XNOR2_X1_LVT multiplier_0i_32_284 (.A(multiplier_0_n_32_89),.B(multiplier_0_n_32_73),.ZN(multiplier_0_n_32_295));
	XNOR2_X1_LVT multiplier_0i_32_285 (.A(multiplier_0_n_32_295),.B(multiplier_0_n_32_57),.ZN(multiplier_0_n_32_296));
	INV_X1_LVT multiplier_0i_32_286 (.A(multiplier_0_n_32_296),.ZN(multiplier_0_n_32_297));
	FA_X1_LVT multiplier_0i_32_299 (.A(multiplier_0_n_32_276),.B(multiplier_0_n_32_304),.CI(multiplier_0_n_32_297),.CO(multiplier_0_n_32_312),.S(multiplier_0_n_32_311));
	FA_X1_LVT multiplier_0i_32_326 (.A(multiplier_0_n_32_318),.B(multiplier_0_n_32_339),.CI(multiplier_0_n_32_312),.CO(multiplier_0_n_32_344),.S(multiplier_0_n_32_343));
	FA_X1_LVT multiplier_0i_32_353 (.A(multiplier_0_n_32_344),.B(multiplier_0_n_32_371),.CI(multiplier_0_n_32_373),.CO(multiplier_0_n_32_376),.S(multiplier_0_n_32_375));
	XNOR2_X1_LVT multiplier_0i_32_276 (.A(multiplier_0_n_32_137),.B(multiplier_0_n_32_121),.ZN(multiplier_0_n_32_287));
	XNOR2_X1_LVT multiplier_0i_32_277 (.A(multiplier_0_n_32_287),.B(multiplier_0_n_32_105),.ZN(multiplier_0_n_32_288));
	OR2_X1_LVT multiplier_0i_32_239 (.A1(multiplier_0_n_32_7),.A2(multiplier_0_n_32_23),.ZN(multiplier_0_n_32_244));
	INV_X1_LVT multiplier_0i_32_241 (.A(multiplier_0_n_32_23),.ZN(multiplier_0_n_32_246));
	NAND2_X1_LVT multiplier_0i_32_240 (.A1(multiplier_0_n_32_211),.A2(multiplier_0_n_32_246),.ZN(multiplier_0_n_32_245));
	INV_X1_LVT multiplier_0i_32_243 (.A(multiplier_0_n_32_7),.ZN(multiplier_0_n_32_248));
	NAND2_X1_LVT multiplier_0i_32_242 (.A1(multiplier_0_n_32_211),.A2(multiplier_0_n_32_248),.ZN(multiplier_0_n_32_247));
	NAND3_X1_LVT multiplier_0i_32_238 (.A1(multiplier_0_n_32_244),.A2(multiplier_0_n_32_245),.A3(multiplier_0_n_32_247),.ZN(multiplier_0_n_32_243));
	XNOR2_X1_LVT multiplier_0i_32_258 (.A(multiplier_0_n_32_56),.B(multiplier_0_n_32_40),.ZN(multiplier_0_n_32_266));
	XNOR2_X1_LVT multiplier_0i_32_259 (.A(multiplier_0_n_32_266),.B(multiplier_0_n_32_24),.ZN(multiplier_0_n_32_267));
	INV_X1_LVT multiplier_0i_32_260 (.A(multiplier_0_n_32_267),.ZN(multiplier_0_n_32_268));
	XNOR2_X1_LVT multiplier_0i_32_251 (.A(multiplier_0_n_32_104),.B(multiplier_0_n_32_88),.ZN(multiplier_0_n_32_259));
	XNOR2_X1_LVT multiplier_0i_32_252 (.A(multiplier_0_n_32_259),.B(multiplier_0_n_32_72),.ZN(multiplier_0_n_32_260));
	INV_X1_LVT multiplier_0i_32_253 (.A(multiplier_0_n_32_260),.ZN(multiplier_0_n_32_261));
	FA_X1_LVT multiplier_0i_32_273 (.A(multiplier_0_n_32_243),.B(multiplier_0_n_32_268),.CI(multiplier_0_n_32_261),.CO(multiplier_0_n_32_282),.S(multiplier_0_n_32_281));
	FA_X1_LVT multiplier_0i_32_300 (.A(multiplier_0_n_32_288),.B(multiplier_0_n_32_309),.CI(multiplier_0_n_32_282),.CO(multiplier_0_n_32_314),.S(multiplier_0_n_32_313));
	FA_X1_LVT multiplier_0i_32_327 (.A(multiplier_0_n_32_314),.B(multiplier_0_n_32_341),.CI(multiplier_0_n_32_343),.CO(multiplier_0_n_32_346),.S(multiplier_0_n_32_345));
	XNOR2_X1_LVT multiplier_0i_32_247 (.A(multiplier_0_n_32_136),.B(multiplier_0_n_32_120),.ZN(multiplier_0_n_32_255));
	INV_X1_LVT multiplier_0i_32_248 (.A(multiplier_0_n_32_255),.ZN(multiplier_0_n_32_256));
	XNOR2_X1_LVT multiplier_0i_32_265 (.A(multiplier_0_n_32_8),.B(multiplier_0_n_32_237),.ZN(multiplier_0_n_32_273));
	XNOR2_X1_LVT multiplier_0i_32_266 (.A(multiplier_0_n_32_273),.B(multiplier_0_n_32_230),.ZN(multiplier_0_n_32_274));
	INV_X1_LVT multiplier_0i_32_267 (.A(multiplier_0_n_32_274),.ZN(multiplier_0_n_32_275));
	FA_X1_LVT multiplier_0i_32_274 (.A(multiplier_0_n_32_256),.B(multiplier_0_n_32_275),.CI(multiplier_0_n_32_250),.CO(multiplier_0_n_32_284),.S(multiplier_0_n_32_283));
	FA_X1_LVT multiplier_0i_32_301 (.A(multiplier_0_n_32_284),.B(multiplier_0_n_32_311),.CI(multiplier_0_n_32_313),.CO(multiplier_0_n_32_316),.S(multiplier_0_n_32_315));
	FA_X1_LVT multiplier_0i_32_275 (.A(multiplier_0_n_32_254),.B(multiplier_0_n_32_252),.CI(multiplier_0_n_32_281),.CO(multiplier_0_n_32_286),.S(multiplier_0_n_32_285));
	FA_X1_LVT multiplier_0i_32_602 (.A(multiplier_0_n_32_283),.B(multiplier_0_n_32_285),.CI(multiplier_0_n_32_658),.CO(multiplier_0_n_32_659),.S(multiplier_0_n_50));
	FA_X1_LVT multiplier_0i_32_603 (.A(multiplier_0_n_32_286),.B(multiplier_0_n_32_315),.CI(multiplier_0_n_32_659),.CO(multiplier_0_n_32_660),.S(multiplier_0_n_51));
	FA_X1_LVT multiplier_0i_32_604 (.A(multiplier_0_n_32_316),.B(multiplier_0_n_32_345),.CI(multiplier_0_n_32_660),.CO(multiplier_0_n_32_661),.S(multiplier_0_n_52));
	FA_X1_LVT multiplier_0i_32_605 (.A(multiplier_0_n_32_346),.B(multiplier_0_n_32_375),.CI(multiplier_0_n_32_661),.CO(multiplier_0_n_32_662),.S(multiplier_0_n_53));
	FA_X1_LVT multiplier_0i_32_606 (.A(multiplier_0_n_32_376),.B(multiplier_0_n_32_405),.CI(multiplier_0_n_32_662),.CO(multiplier_0_n_32_663),.S(multiplier_0_n_54));
	FA_X1_LVT multiplier_0i_32_607 (.A(multiplier_0_n_32_406),.B(multiplier_0_n_32_435),.CI(multiplier_0_n_32_663),.CO(multiplier_0_n_32_664),.S(multiplier_0_n_55));
	FA_X1_LVT multiplier_0i_32_608 (.A(multiplier_0_n_32_436),.B(multiplier_0_n_32_465),.CI(multiplier_0_n_32_664),.CO(multiplier_0_n_32_665),.S(multiplier_0_n_56));
	FA_X1_LVT multiplier_0i_32_609 (.A(multiplier_0_n_32_466),.B(multiplier_0_n_32_495),.CI(multiplier_0_n_32_665),.CO(multiplier_0_n_32_666),.S(multiplier_0_n_57));
	INV_X1_LVT multiplier_0i_34_31 (.A(multiplier_0_n_57),.ZN(multiplier_0_n_34_16));
	OAI22_X1_LVT multiplier_0i_34_32 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_7),.B1(multiplier_0_n_34_16),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[15]));
	INV_X1_LVT multiplier_0i_34_12 (.A(multiplier_0_n_48),.ZN(multiplier_0_n_34_6));
	INV_X1_LVT multiplier_0i_34_29 (.A(multiplier_0_n_56),.ZN(multiplier_0_n_34_15));
	OAI22_X1_LVT multiplier_0i_34_30 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_6),.B1(multiplier_0_n_34_15),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[14]));
	AOI22_X1_LVT multiplier_0i_45_29 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_136),.B1(multiplier_0_reslo_wr),.B2(multiplier_0_per_din_msk[14]),.ZN(multiplier_0_n_45_15));
	INV_X1_LVT multiplier_0i_45_30 (.A(multiplier_0_n_45_15),.ZN(multiplier_0_n_119));
	OR2_X1_LVT multiplier_0i_23_0 (.A1(multiplier_0_cycle[0]),.A2(multiplier_0_cycle[1]),.ZN(multiplier_0_result_wr));
	INV_X1_LVT multiplier_0i_39_1 (.A(multiplier_0_result_wr),.ZN(multiplier_0_n_39_1));
	INV_X1_LVT multiplier_0i_39_0 (.A(multiplier_0_result_clr),.ZN(multiplier_0_n_39_0));
	NAND2_X1_LVT multiplier_0i_39_2 (.A1(multiplier_0_n_39_1),.A2(multiplier_0_n_39_0),.ZN(multiplier_0_n_69));
	INV_X1_LVT multiplier_0i_46_1 (.A(multiplier_0_n_69),.ZN(multiplier_0_n_46_1));
	INV_X1_LVT multiplier_0i_46_0 (.A(multiplier_0_reslo_wr),.ZN(multiplier_0_n_46_0));
	NAND2_X1_LVT multiplier_0i_46_2 (.A1(multiplier_0_n_46_1),.A2(multiplier_0_n_46_0),.ZN(multiplier_0_n_121));
	CLKGATETST_X1_LVT multiplier_0clk_gate_reslo_reg (.CK(mclk),.E(multiplier_0_n_121),.SE(1'b0),.GCK(multiplier_0_n_88));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b14___05F05d (.D(multiplier_0_n_119),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_90),.QN());
	INV_X1_LVT multiplier_0i_34_10 (.A(multiplier_0_n_47),.ZN(multiplier_0_n_34_5));
	INV_X1_LVT multiplier_0i_34_27 (.A(multiplier_0_n_55),.ZN(multiplier_0_n_34_14));
	OAI22_X1_LVT multiplier_0i_34_28 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_5),.B1(multiplier_0_n_34_14),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[13]));
	AOI22_X1_LVT multiplier_0i_45_27 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_135),.B1(multiplier_0_reslo_wr),.B2(multiplier_0_per_din_msk[13]),.ZN(multiplier_0_n_45_14));
	INV_X1_LVT multiplier_0i_45_28 (.A(multiplier_0_n_45_14),.ZN(multiplier_0_n_118));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b13___05F05d (.D(multiplier_0_n_118),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_91),.QN());
	INV_X1_LVT multiplier_0i_34_8 (.A(multiplier_0_n_46),.ZN(multiplier_0_n_34_4));
	INV_X1_LVT multiplier_0i_34_25 (.A(multiplier_0_n_54),.ZN(multiplier_0_n_34_13));
	OAI22_X1_LVT multiplier_0i_34_26 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_4),.B1(multiplier_0_n_34_13),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[12]));
	AOI22_X1_LVT multiplier_0i_45_25 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_134),.B1(multiplier_0_reslo_wr),.B2(multiplier_0_per_din_msk[12]),.ZN(multiplier_0_n_45_13));
	INV_X1_LVT multiplier_0i_45_26 (.A(multiplier_0_n_45_13),.ZN(multiplier_0_n_117));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b12___05F05d (.D(multiplier_0_n_117),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_92),.QN());
	INV_X1_LVT multiplier_0i_34_6 (.A(multiplier_0_n_45),.ZN(multiplier_0_n_34_3));
	INV_X1_LVT multiplier_0i_34_23 (.A(multiplier_0_n_53),.ZN(multiplier_0_n_34_12));
	OAI22_X1_LVT multiplier_0i_34_24 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_3),.B1(multiplier_0_n_34_12),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[11]));
	AOI22_X1_LVT multiplier_0i_45_23 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_133),.B1(multiplier_0_reslo_wr),.B2(multiplier_0_per_din_msk[11]),.ZN(multiplier_0_n_45_12));
	INV_X1_LVT multiplier_0i_45_24 (.A(multiplier_0_n_45_12),.ZN(multiplier_0_n_116));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b11___05F05d (.D(multiplier_0_n_116),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_93),.QN());
	XNOR2_X1_LVT multiplier_0i_32_589 (.A(multiplier_0_n_32_2),.B(multiplier_0_n_32_153),.ZN(multiplier_0_n_32_647));
	XNOR2_X1_LVT multiplier_0i_32_590 (.A(multiplier_0_n_32_647),.B(multiplier_0_n_32_646),.ZN(multiplier_0_n_32_648));
	INV_X1_LVT multiplier_0i_32_591 (.A(multiplier_0_n_32_648),.ZN(multiplier_0_n_44));
	INV_X1_LVT multiplier_0i_34_4 (.A(multiplier_0_n_44),.ZN(multiplier_0_n_34_2));
	INV_X1_LVT multiplier_0i_34_21 (.A(multiplier_0_n_52),.ZN(multiplier_0_n_34_11));
	OAI22_X1_LVT multiplier_0i_34_22 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_2),.B1(multiplier_0_n_34_11),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[10]));
	AOI22_X1_LVT multiplier_0i_45_21 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_132),.B1(multiplier_0_reslo_wr),.B2(multiplier_0_per_din_msk[10]),.ZN(multiplier_0_n_45_11));
	INV_X1_LVT multiplier_0i_45_22 (.A(multiplier_0_n_45_11),.ZN(multiplier_0_n_115));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b10___05F05d (.D(multiplier_0_n_115),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_94),.QN());
	XNOR2_X1_LVT multiplier_0i_32_586 (.A(multiplier_0_n_32_17),.B(multiplier_0_n_32_1),.ZN(multiplier_0_n_32_645));
	INV_X1_LVT multiplier_0i_32_587 (.A(multiplier_0_n_32_645),.ZN(multiplier_0_n_43));
	INV_X1_LVT multiplier_0i_34_2 (.A(multiplier_0_n_43),.ZN(multiplier_0_n_34_1));
	INV_X1_LVT multiplier_0i_34_19 (.A(multiplier_0_n_51),.ZN(multiplier_0_n_34_10));
	OAI22_X1_LVT multiplier_0i_34_20 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_1),.B1(multiplier_0_n_34_10),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[9]));
	AOI22_X1_LVT multiplier_0i_45_19 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_131),.B1(multiplier_0_reslo_wr),.B2(multiplier_0_per_din_msk[9]),.ZN(multiplier_0_n_45_10));
	INV_X1_LVT multiplier_0i_45_20 (.A(multiplier_0_n_45_10),.ZN(multiplier_0_n_114));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b9___05F05d (.D(multiplier_0_n_114),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_95),.QN());
	NAND2_X1_LVT multiplier_0i_32_0 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1[0]),.ZN(multiplier_0_n_32_0));
	INV_X1_LVT multiplier_0i_32_585 (.A(multiplier_0_n_32_0),.ZN(multiplier_0_n_42));
	INV_X1_LVT multiplier_0i_34_0 (.A(multiplier_0_n_42),.ZN(multiplier_0_n_34_0));
	INV_X1_LVT multiplier_0i_34_17 (.A(multiplier_0_n_50),.ZN(multiplier_0_n_34_9));
	OAI22_X1_LVT multiplier_0i_34_18 (.A1(multiplier_0_n_34_0),.A2(multiplier_0_n_34_8),.B1(multiplier_0_n_34_9),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[8]));
	AOI22_X1_LVT multiplier_0i_45_17 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_130),.B1(multiplier_0_reslo_wr),.B2(multiplier_0_per_din_msk[8]),.ZN(multiplier_0_n_45_9));
	INV_X1_LVT multiplier_0i_45_18 (.A(multiplier_0_n_45_9),.ZN(multiplier_0_n_113));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b8___05F05d (.D(multiplier_0_n_113),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_96),.QN());
	NOR2_X1_LVT multiplier_0i_34_15 (.A1(multiplier_0_n_34_7),.A2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[7]));
	AOI22_X1_LVT multiplier_0i_45_15 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_129),.B1(multiplier_0_reslo_wr),.B2(per_din[7]),.ZN(multiplier_0_n_45_8));
	INV_X1_LVT multiplier_0i_45_16 (.A(multiplier_0_n_45_8),.ZN(multiplier_0_n_112));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b7___05F05d (.D(multiplier_0_n_112),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_97),.QN());
	NOR2_X1_LVT multiplier_0i_34_13 (.A1(multiplier_0_n_34_6),.A2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[6]));
	AOI22_X1_LVT multiplier_0i_45_13 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_128),.B1(multiplier_0_reslo_wr),.B2(per_din[6]),.ZN(multiplier_0_n_45_7));
	INV_X1_LVT multiplier_0i_45_14 (.A(multiplier_0_n_45_7),.ZN(multiplier_0_n_111));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b6___05F05d (.D(multiplier_0_n_111),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_98),.QN());
	NOR2_X1_LVT multiplier_0i_34_11 (.A1(multiplier_0_n_34_5),.A2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[5]));
	AOI22_X1_LVT multiplier_0i_45_11 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_127),.B1(multiplier_0_reslo_wr),.B2(per_din[5]),.ZN(multiplier_0_n_45_6));
	INV_X1_LVT multiplier_0i_45_12 (.A(multiplier_0_n_45_6),.ZN(multiplier_0_n_110));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b5___05F05d (.D(multiplier_0_n_110),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_99),.QN());
	NOR2_X1_LVT multiplier_0i_34_9 (.A1(multiplier_0_n_34_4),.A2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[4]));
	AOI22_X1_LVT multiplier_0i_45_9 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_126),.B1(multiplier_0_reslo_wr),.B2(per_din[4]),.ZN(multiplier_0_n_45_5));
	INV_X1_LVT multiplier_0i_45_10 (.A(multiplier_0_n_45_5),.ZN(multiplier_0_n_109));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b4___05F05d (.D(multiplier_0_n_109),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_100),.QN());
	NOR2_X1_LVT multiplier_0i_34_7 (.A1(multiplier_0_n_34_3),.A2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[3]));
	AOI22_X1_LVT multiplier_0i_45_7 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_125),.B1(multiplier_0_reslo_wr),.B2(per_din[3]),.ZN(multiplier_0_n_45_4));
	INV_X1_LVT multiplier_0i_45_8 (.A(multiplier_0_n_45_4),.ZN(multiplier_0_n_108));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b3___05F05d (.D(multiplier_0_n_108),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_101),.QN());
	NOR2_X1_LVT multiplier_0i_34_5 (.A1(multiplier_0_n_34_2),.A2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[2]));
	AOI22_X1_LVT multiplier_0i_45_5 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_124),.B1(multiplier_0_reslo_wr),.B2(per_din[2]),.ZN(multiplier_0_n_45_3));
	INV_X1_LVT multiplier_0i_45_6 (.A(multiplier_0_n_45_3),.ZN(multiplier_0_n_107));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b2___05F05d (.D(multiplier_0_n_107),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_102),.QN());
	NOR2_X1_LVT multiplier_0i_34_3 (.A1(multiplier_0_n_34_1),.A2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[1]));
	AOI22_X1_LVT multiplier_0i_45_3 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_123),.B1(multiplier_0_reslo_wr),.B2(per_din[1]),.ZN(multiplier_0_n_45_2));
	INV_X1_LVT multiplier_0i_45_4 (.A(multiplier_0_n_45_2),.ZN(multiplier_0_n_106));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b1___05F05d (.D(multiplier_0_n_106),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_103),.QN());
	NOR2_X1_LVT multiplier_0i_34_1 (.A1(multiplier_0_n_34_0),.A2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_45_1 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_122),.B1(per_din[0]),.B2(multiplier_0_reslo_wr),.ZN(multiplier_0_n_45_1));
	INV_X1_LVT multiplier_0i_45_2 (.A(multiplier_0_n_45_1),.ZN(multiplier_0_n_105));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b0___05F05d (.D(multiplier_0_n_105),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_104),.QN());
	HA_X1_LVT multiplier_0i_48_0 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_n_104),.CO(multiplier_0_n_48_0),.S(multiplier_0_n_122));
	FA_X1_LVT multiplier_0i_48_1 (.A(multiplier_0_product_xp[1]),.B(multiplier_0_n_103),.CI(multiplier_0_n_48_0),.CO(multiplier_0_n_48_1),.S(multiplier_0_n_123));
	FA_X1_LVT multiplier_0i_48_2 (.A(multiplier_0_product_xp[2]),.B(multiplier_0_n_102),.CI(multiplier_0_n_48_1),.CO(multiplier_0_n_48_2),.S(multiplier_0_n_124));
	FA_X1_LVT multiplier_0i_48_3 (.A(multiplier_0_product_xp[3]),.B(multiplier_0_n_101),.CI(multiplier_0_n_48_2),.CO(multiplier_0_n_48_3),.S(multiplier_0_n_125));
	FA_X1_LVT multiplier_0i_48_4 (.A(multiplier_0_product_xp[4]),.B(multiplier_0_n_100),.CI(multiplier_0_n_48_3),.CO(multiplier_0_n_48_4),.S(multiplier_0_n_126));
	FA_X1_LVT multiplier_0i_48_5 (.A(multiplier_0_product_xp[5]),.B(multiplier_0_n_99),.CI(multiplier_0_n_48_4),.CO(multiplier_0_n_48_5),.S(multiplier_0_n_127));
	FA_X1_LVT multiplier_0i_48_6 (.A(multiplier_0_product_xp[6]),.B(multiplier_0_n_98),.CI(multiplier_0_n_48_5),.CO(multiplier_0_n_48_6),.S(multiplier_0_n_128));
	FA_X1_LVT multiplier_0i_48_7 (.A(multiplier_0_product_xp[7]),.B(multiplier_0_n_97),.CI(multiplier_0_n_48_6),.CO(multiplier_0_n_48_7),.S(multiplier_0_n_129));
	FA_X1_LVT multiplier_0i_48_8 (.A(multiplier_0_product_xp[8]),.B(multiplier_0_n_96),.CI(multiplier_0_n_48_7),.CO(multiplier_0_n_48_8),.S(multiplier_0_n_130));
	FA_X1_LVT multiplier_0i_48_9 (.A(multiplier_0_product_xp[9]),.B(multiplier_0_n_95),.CI(multiplier_0_n_48_8),.CO(multiplier_0_n_48_9),.S(multiplier_0_n_131));
	FA_X1_LVT multiplier_0i_48_10 (.A(multiplier_0_product_xp[10]),.B(multiplier_0_n_94),.CI(multiplier_0_n_48_9),.CO(multiplier_0_n_48_10),.S(multiplier_0_n_132));
	FA_X1_LVT multiplier_0i_48_11 (.A(multiplier_0_product_xp[11]),.B(multiplier_0_n_93),.CI(multiplier_0_n_48_10),.CO(multiplier_0_n_48_11),.S(multiplier_0_n_133));
	FA_X1_LVT multiplier_0i_48_12 (.A(multiplier_0_product_xp[12]),.B(multiplier_0_n_92),.CI(multiplier_0_n_48_11),.CO(multiplier_0_n_48_12),.S(multiplier_0_n_134));
	FA_X1_LVT multiplier_0i_48_13 (.A(multiplier_0_product_xp[13]),.B(multiplier_0_n_91),.CI(multiplier_0_n_48_12),.CO(multiplier_0_n_48_13),.S(multiplier_0_n_135));
	FA_X1_LVT multiplier_0i_48_14 (.A(multiplier_0_product_xp[14]),.B(multiplier_0_n_90),.CI(multiplier_0_n_48_13),.CO(multiplier_0_n_48_14),.S(multiplier_0_n_136));
	FA_X1_LVT multiplier_0i_48_15 (.A(multiplier_0_product_xp[15]),.B(multiplier_0_n_89),.CI(multiplier_0_n_48_14),.CO(multiplier_0_n_48_15),.S(multiplier_0_n_137));
	AOI22_X1_LVT multiplier_0i_45_31 (.A1(multiplier_0_n_45_0),.A2(multiplier_0_n_137),.B1(multiplier_0_reslo_wr),.B2(multiplier_0_per_din_msk[15]),.ZN(multiplier_0_n_45_16));
	INV_X1_LVT multiplier_0i_45_32 (.A(multiplier_0_n_45_16),.ZN(multiplier_0_n_120));
	DFFR_X1_LVT multiplier_0reslo_reg___05F05b15___05F05d (.D(multiplier_0_n_120),.RN(multiplier_0_n_38),.CK(multiplier_0_n_88),.Q(multiplier_0_n_89),.QN());
	AOI22_X1_LVT multiplier_0i_60_93 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_89),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_137),.ZN(multiplier_0_n_60_78));
	NOR2_X1_LVT multiplier_0i_1_0 (.A1(per_we[0]),.A2(per_we[1]),.ZN(multiplier_0_n_0));
	AND2_X1_LVT multiplier_0i_2_0 (.A1(multiplier_0_n_0),.A2(multiplier_0_reg_sel),.ZN(multiplier_0_reg_read));
	AND2_X1_LVT multiplier_0i_4_5 (.A1(multiplier_0_reg_read),.A2(multiplier_0_n_6),.ZN(multiplier_0_n_13));
	INV_X1_LVT multiplier_0i_60_2 (.A(multiplier_0_n_13),.ZN(multiplier_0_n_60_2));
	NOR2_X1_LVT multiplier_0i_60_94 (.A1(multiplier_0_n_60_78),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_79));
	AND2_X1_LVT multiplier_0i_4_0 (.A1(multiplier_0_n_1),.A2(multiplier_0_reg_read),.ZN(multiplier_0_n_9));
	AND2_X1_LVT multiplier_0i_4_3 (.A1(multiplier_0_reg_read),.A2(multiplier_0_n_4),.ZN(multiplier_0_n_11));
	AND2_X1_LVT multiplier_0i_4_2 (.A1(multiplier_0_reg_read),.A2(multiplier_0_n_3),.ZN(multiplier_0_reg_rd1));
	AND2_X1_LVT multiplier_0i_4_1 (.A1(multiplier_0_reg_read),.A2(multiplier_0_n_2),.ZN(multiplier_0_n_10));
	OR4_X1_LVT multiplier_0i_59_0 (.A1(multiplier_0_n_9),.A2(multiplier_0_n_11),.A3(multiplier_0_reg_rd1),.A4(multiplier_0_n_10),.ZN(multiplier_0_n_150));
	AND2_X1_LVT multiplier_0i_60_95 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_60_80));
	INV_X1_LVT multiplier_0i_57_0 (.A(multiplier_0_cycle[1]),.ZN(multiplier_0_n_57_0));
	INV_X1_LVT multiplier_0i_52_0 (.A(multiplier_0_op2_wr),.ZN(multiplier_0_n_52_0));
	NAND2_X1_LVT multiplier_0i_32_151 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_32_151));
	AND2_X1_LVT multiplier_0i_31_0 (.A1(multiplier_0_op1[15]),.A2(multiplier_0_sign_sel),.ZN(multiplier_0_op1_xp[0]));
	NAND2_X1_LVT multiplier_0i_32_135 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1_xp[0]),.ZN(multiplier_0_n_32_135));
	XNOR2_X1_LVT multiplier_0i_32_583 (.A(multiplier_0_n_32_151),.B(multiplier_0_n_32_135),.ZN(multiplier_0_n_32_643));
	NAND2_X1_LVT multiplier_0i_32_150 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_32_150));
	NAND2_X1_LVT multiplier_0i_32_134 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_32_134));
	INV_X1_LVT multiplier_0i_32_579 (.A(multiplier_0_n_32_134),.ZN(multiplier_0_n_32_638));
	NAND2_X1_LVT multiplier_0i_32_578 (.A1(multiplier_0_n_32_150),.A2(multiplier_0_n_32_638),.ZN(multiplier_0_n_32_637));
	NAND2_X1_LVT multiplier_0i_32_118 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1_xp[0]),.ZN(multiplier_0_n_32_118));
	NAND2_X1_LVT multiplier_0i_32_580 (.A1(multiplier_0_n_32_118),.A2(multiplier_0_n_32_150),.ZN(multiplier_0_n_32_639));
	NAND2_X1_LVT multiplier_0i_32_581 (.A1(multiplier_0_n_32_118),.A2(multiplier_0_n_32_638),.ZN(multiplier_0_n_32_640));
	NAND3_X1_LVT multiplier_0i_32_577 (.A1(multiplier_0_n_32_637),.A2(multiplier_0_n_32_639),.A3(multiplier_0_n_32_640),.ZN(multiplier_0_n_32_636));
	XNOR2_X1_LVT multiplier_0i_32_584 (.A(multiplier_0_n_32_643),.B(multiplier_0_n_32_636),.ZN(multiplier_0_n_32_644));
	NAND2_X1_LVT multiplier_0i_32_149 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_32_149));
	NAND2_X1_LVT multiplier_0i_32_133 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_32_133));
	INV_X1_LVT multiplier_0i_32_568 (.A(multiplier_0_n_32_133),.ZN(multiplier_0_n_32_625));
	NAND2_X1_LVT multiplier_0i_32_567 (.A1(multiplier_0_n_32_149),.A2(multiplier_0_n_32_625),.ZN(multiplier_0_n_32_624));
	NAND2_X1_LVT multiplier_0i_32_117 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_32_117));
	INV_X1_LVT multiplier_0i_32_570 (.A(multiplier_0_n_32_117),.ZN(multiplier_0_n_32_627));
	NAND2_X1_LVT multiplier_0i_32_569 (.A1(multiplier_0_n_32_149),.A2(multiplier_0_n_32_627),.ZN(multiplier_0_n_32_626));
	OR2_X1_LVT multiplier_0i_32_571 (.A1(multiplier_0_n_32_117),.A2(multiplier_0_n_32_133),.ZN(multiplier_0_n_32_628));
	NAND3_X1_LVT multiplier_0i_32_566 (.A1(multiplier_0_n_32_624),.A2(multiplier_0_n_32_626),.A3(multiplier_0_n_32_628),.ZN(multiplier_0_n_32_623));
	NAND2_X1_LVT multiplier_0i_32_101 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1_xp[0]),.ZN(multiplier_0_n_32_101));
	NAND2_X1_LVT multiplier_0i_32_148 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_32_148));
	NAND2_X1_LVT multiplier_0i_32_132 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_32_132));
	INV_X1_LVT multiplier_0i_32_550 (.A(multiplier_0_n_32_132),.ZN(multiplier_0_n_32_605));
	NAND2_X1_LVT multiplier_0i_32_549 (.A1(multiplier_0_n_32_148),.A2(multiplier_0_n_32_605),.ZN(multiplier_0_n_32_604));
	NAND2_X1_LVT multiplier_0i_32_116 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_32_116));
	INV_X1_LVT multiplier_0i_32_552 (.A(multiplier_0_n_32_116),.ZN(multiplier_0_n_32_607));
	NAND2_X1_LVT multiplier_0i_32_551 (.A1(multiplier_0_n_32_148),.A2(multiplier_0_n_32_607),.ZN(multiplier_0_n_32_606));
	OR2_X1_LVT multiplier_0i_32_553 (.A1(multiplier_0_n_32_116),.A2(multiplier_0_n_32_132),.ZN(multiplier_0_n_32_608));
	NAND3_X1_LVT multiplier_0i_32_548 (.A1(multiplier_0_n_32_604),.A2(multiplier_0_n_32_606),.A3(multiplier_0_n_32_608),.ZN(multiplier_0_n_32_603));
	NAND2_X1_LVT multiplier_0i_32_84 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1_xp[0]),.ZN(multiplier_0_n_32_84));
	NAND2_X1_LVT multiplier_0i_32_100 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_32_100));
	INV_X1_LVT multiplier_0i_32_559 (.A(multiplier_0_n_32_100),.ZN(multiplier_0_n_32_614));
	NAND2_X1_LVT multiplier_0i_32_558 (.A1(multiplier_0_n_32_84),.A2(multiplier_0_n_32_614),.ZN(multiplier_0_n_32_613));
	NAND2_X1_LVT multiplier_0i_32_83 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_32_83));
	NAND2_X1_LVT multiplier_0i_32_99 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_32_99));
	OR2_X1_LVT multiplier_0i_32_538 (.A1(multiplier_0_n_32_83),.A2(multiplier_0_n_32_99),.ZN(multiplier_0_n_32_590));
	NAND2_X1_LVT multiplier_0i_32_67 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1_xp[0]),.ZN(multiplier_0_n_32_67));
	INV_X1_LVT multiplier_0i_32_540 (.A(multiplier_0_n_32_99),.ZN(multiplier_0_n_32_592));
	NAND2_X1_LVT multiplier_0i_32_539 (.A1(multiplier_0_n_32_67),.A2(multiplier_0_n_32_592),.ZN(multiplier_0_n_32_591));
	INV_X1_LVT multiplier_0i_32_542 (.A(multiplier_0_n_32_83),.ZN(multiplier_0_n_32_594));
	NAND2_X1_LVT multiplier_0i_32_541 (.A1(multiplier_0_n_32_67),.A2(multiplier_0_n_32_594),.ZN(multiplier_0_n_32_593));
	NAND3_X1_LVT multiplier_0i_32_537 (.A1(multiplier_0_n_32_590),.A2(multiplier_0_n_32_591),.A3(multiplier_0_n_32_593),.ZN(multiplier_0_n_32_589));
	NAND2_X1_LVT multiplier_0i_32_560 (.A1(multiplier_0_n_32_589),.A2(multiplier_0_n_32_614),.ZN(multiplier_0_n_32_615));
	NAND2_X1_LVT multiplier_0i_32_561 (.A1(multiplier_0_n_32_589),.A2(multiplier_0_n_32_84),.ZN(multiplier_0_n_32_616));
	NAND3_X1_LVT multiplier_0i_32_557 (.A1(multiplier_0_n_32_613),.A2(multiplier_0_n_32_615),.A3(multiplier_0_n_32_616),.ZN(multiplier_0_n_32_612));
	FA_X1_LVT multiplier_0i_32_572 (.A(multiplier_0_n_32_101),.B(multiplier_0_n_32_603),.CI(multiplier_0_n_32_612),.CO(multiplier_0_n_32_630),.S(multiplier_0_n_32_629));
	XNOR2_X1_LVT multiplier_0i_32_574 (.A(multiplier_0_n_32_150),.B(multiplier_0_n_32_134),.ZN(multiplier_0_n_32_633));
	XNOR2_X1_LVT multiplier_0i_32_575 (.A(multiplier_0_n_32_633),.B(multiplier_0_n_32_118),.ZN(multiplier_0_n_32_634));
	INV_X1_LVT multiplier_0i_32_576 (.A(multiplier_0_n_32_634),.ZN(multiplier_0_n_32_635));
	FA_X1_LVT multiplier_0i_32_582 (.A(multiplier_0_n_32_623),.B(multiplier_0_n_32_630),.CI(multiplier_0_n_32_635),.CO(multiplier_0_n_32_642),.S(multiplier_0_n_32_641));
	XNOR2_X1_LVT multiplier_0i_32_617 (.A(multiplier_0_n_32_644),.B(multiplier_0_n_32_642),.ZN(multiplier_0_n_32_674));
	XNOR2_X1_LVT multiplier_0i_32_564 (.A(multiplier_0_n_32_149),.B(multiplier_0_n_32_133),.ZN(multiplier_0_n_32_621));
	XNOR2_X1_LVT multiplier_0i_32_565 (.A(multiplier_0_n_32_621),.B(multiplier_0_n_32_117),.ZN(multiplier_0_n_32_622));
	NAND2_X1_LVT multiplier_0i_32_147 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_32_147));
	NAND2_X1_LVT multiplier_0i_32_131 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_32_131));
	INV_X1_LVT multiplier_0i_32_531 (.A(multiplier_0_n_32_131),.ZN(multiplier_0_n_32_583));
	NAND2_X1_LVT multiplier_0i_32_530 (.A1(multiplier_0_n_32_147),.A2(multiplier_0_n_32_583),.ZN(multiplier_0_n_32_582));
	NAND2_X1_LVT multiplier_0i_32_115 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_32_115));
	INV_X1_LVT multiplier_0i_32_533 (.A(multiplier_0_n_32_115),.ZN(multiplier_0_n_32_585));
	NAND2_X1_LVT multiplier_0i_32_532 (.A1(multiplier_0_n_32_147),.A2(multiplier_0_n_32_585),.ZN(multiplier_0_n_32_584));
	OR2_X1_LVT multiplier_0i_32_534 (.A1(multiplier_0_n_32_115),.A2(multiplier_0_n_32_131),.ZN(multiplier_0_n_32_586));
	NAND3_X1_LVT multiplier_0i_32_529 (.A1(multiplier_0_n_32_582),.A2(multiplier_0_n_32_584),.A3(multiplier_0_n_32_586),.ZN(multiplier_0_n_32_581));
	NAND2_X1_LVT multiplier_0i_32_82 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_32_82));
	NAND2_X1_LVT multiplier_0i_32_98 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_32_98));
	NOR2_X1_LVT multiplier_0i_32_520 (.A1(multiplier_0_n_32_82),.A2(multiplier_0_n_32_98),.ZN(multiplier_0_n_32_568));
	NAND2_X1_LVT multiplier_0i_32_66 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_32_66));
	NOR2_X1_LVT multiplier_0i_32_521 (.A1(multiplier_0_n_32_66),.A2(multiplier_0_n_32_98),.ZN(multiplier_0_n_32_569));
	NOR2_X1_LVT multiplier_0i_32_522 (.A1(multiplier_0_n_32_66),.A2(multiplier_0_n_32_82),.ZN(multiplier_0_n_32_570));
	OR3_X1_LVT multiplier_0i_32_519 (.A1(multiplier_0_n_32_568),.A2(multiplier_0_n_32_569),.A3(multiplier_0_n_32_570),.ZN(multiplier_0_n_32_567));
	NAND2_X1_LVT multiplier_0i_32_146 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_32_146));
	NAND2_X1_LVT multiplier_0i_32_130 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_32_130));
	INV_X1_LVT multiplier_0i_32_512 (.A(multiplier_0_n_32_130),.ZN(multiplier_0_n_32_560));
	NAND2_X1_LVT multiplier_0i_32_511 (.A1(multiplier_0_n_32_146),.A2(multiplier_0_n_32_560),.ZN(multiplier_0_n_32_559));
	NAND2_X1_LVT multiplier_0i_32_114 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_32_114));
	INV_X1_LVT multiplier_0i_32_514 (.A(multiplier_0_n_32_114),.ZN(multiplier_0_n_32_562));
	NAND2_X1_LVT multiplier_0i_32_513 (.A1(multiplier_0_n_32_146),.A2(multiplier_0_n_32_562),.ZN(multiplier_0_n_32_561));
	OR2_X1_LVT multiplier_0i_32_515 (.A1(multiplier_0_n_32_114),.A2(multiplier_0_n_32_130),.ZN(multiplier_0_n_32_563));
	NAND3_X1_LVT multiplier_0i_32_510 (.A1(multiplier_0_n_32_559),.A2(multiplier_0_n_32_561),.A3(multiplier_0_n_32_563),.ZN(multiplier_0_n_32_558));
	NAND2_X1_LVT multiplier_0i_32_50 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1_xp[0]),.ZN(multiplier_0_n_32_50));
	NAND2_X1_LVT multiplier_0i_32_81 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_32_81));
	NAND2_X1_LVT multiplier_0i_32_97 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_32_97));
	NOR2_X1_LVT multiplier_0i_32_493 (.A1(multiplier_0_n_32_81),.A2(multiplier_0_n_32_97),.ZN(multiplier_0_n_32_537));
	NAND2_X1_LVT multiplier_0i_32_65 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_32_65));
	NOR2_X1_LVT multiplier_0i_32_494 (.A1(multiplier_0_n_32_65),.A2(multiplier_0_n_32_97),.ZN(multiplier_0_n_32_538));
	NOR2_X1_LVT multiplier_0i_32_495 (.A1(multiplier_0_n_32_65),.A2(multiplier_0_n_32_81),.ZN(multiplier_0_n_32_539));
	OR3_X1_LVT multiplier_0i_32_492 (.A1(multiplier_0_n_32_537),.A2(multiplier_0_n_32_538),.A3(multiplier_0_n_32_539),.ZN(multiplier_0_n_32_536));
	NAND2_X1_LVT multiplier_0i_32_145 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_32_145));
	NAND2_X1_LVT multiplier_0i_32_129 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_32_129));
	INV_X1_LVT multiplier_0i_32_485 (.A(multiplier_0_n_32_129),.ZN(multiplier_0_n_32_529));
	NAND2_X1_LVT multiplier_0i_32_484 (.A1(multiplier_0_n_32_145),.A2(multiplier_0_n_32_529),.ZN(multiplier_0_n_32_528));
	NAND2_X1_LVT multiplier_0i_32_113 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_32_113));
	INV_X1_LVT multiplier_0i_32_487 (.A(multiplier_0_n_32_113),.ZN(multiplier_0_n_32_531));
	NAND2_X1_LVT multiplier_0i_32_486 (.A1(multiplier_0_n_32_145),.A2(multiplier_0_n_32_531),.ZN(multiplier_0_n_32_530));
	OR2_X1_LVT multiplier_0i_32_488 (.A1(multiplier_0_n_32_113),.A2(multiplier_0_n_32_129),.ZN(multiplier_0_n_32_532));
	NAND3_X1_LVT multiplier_0i_32_483 (.A1(multiplier_0_n_32_528),.A2(multiplier_0_n_32_530),.A3(multiplier_0_n_32_532),.ZN(multiplier_0_n_32_527));
	FA_X1_LVT multiplier_0i_32_523 (.A(multiplier_0_n_32_50),.B(multiplier_0_n_32_536),.CI(multiplier_0_n_32_527),.CO(multiplier_0_n_32_572),.S(multiplier_0_n_32_571));
	FA_X1_LVT multiplier_0i_32_543 (.A(multiplier_0_n_32_567),.B(multiplier_0_n_32_558),.CI(multiplier_0_n_32_572),.CO(multiplier_0_n_32_596),.S(multiplier_0_n_32_595));
	XNOR2_X1_LVT multiplier_0i_32_554 (.A(multiplier_0_n_32_100),.B(multiplier_0_n_32_84),.ZN(multiplier_0_n_32_609));
	XNOR2_X1_LVT multiplier_0i_32_555 (.A(multiplier_0_n_32_609),.B(multiplier_0_n_32_589),.ZN(multiplier_0_n_32_610));
	INV_X1_LVT multiplier_0i_32_556 (.A(multiplier_0_n_32_610),.ZN(multiplier_0_n_32_611));
	FA_X1_LVT multiplier_0i_32_562 (.A(multiplier_0_n_32_581),.B(multiplier_0_n_32_596),.CI(multiplier_0_n_32_611),.CO(multiplier_0_n_32_618),.S(multiplier_0_n_32_617));
	FA_X1_LVT multiplier_0i_32_573 (.A(multiplier_0_n_32_622),.B(multiplier_0_n_32_629),.CI(multiplier_0_n_32_618),.CO(multiplier_0_n_32_632),.S(multiplier_0_n_32_631));
	XNOR2_X1_LVT multiplier_0i_32_546 (.A(multiplier_0_n_32_148),.B(multiplier_0_n_32_132),.ZN(multiplier_0_n_32_601));
	XNOR2_X1_LVT multiplier_0i_32_547 (.A(multiplier_0_n_32_601),.B(multiplier_0_n_32_116),.ZN(multiplier_0_n_32_602));
	XNOR2_X1_LVT multiplier_0i_32_535 (.A(multiplier_0_n_32_99),.B(multiplier_0_n_32_83),.ZN(multiplier_0_n_32_587));
	XNOR2_X1_LVT multiplier_0i_32_536 (.A(multiplier_0_n_32_587),.B(multiplier_0_n_32_67),.ZN(multiplier_0_n_32_588));
	XNOR2_X1_LVT multiplier_0i_32_527 (.A(multiplier_0_n_32_147),.B(multiplier_0_n_32_131),.ZN(multiplier_0_n_32_579));
	XNOR2_X1_LVT multiplier_0i_32_528 (.A(multiplier_0_n_32_579),.B(multiplier_0_n_32_115),.ZN(multiplier_0_n_32_580));
	FA_X1_LVT multiplier_0i_32_544 (.A(multiplier_0_n_32_588),.B(multiplier_0_n_32_580),.CI(multiplier_0_n_32_595),.CO(multiplier_0_n_32_598),.S(multiplier_0_n_32_597));
	FA_X1_LVT multiplier_0i_32_563 (.A(multiplier_0_n_32_602),.B(multiplier_0_n_32_598),.CI(multiplier_0_n_32_617),.CO(multiplier_0_n_32_620),.S(multiplier_0_n_32_619));
	NAND2_X1_LVT multiplier_0i_32_33 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1_xp[0]),.ZN(multiplier_0_n_32_33));
	NAND2_X1_LVT multiplier_0i_32_49 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_32_49));
	INV_X1_LVT multiplier_0i_32_501 (.A(multiplier_0_n_32_49),.ZN(multiplier_0_n_32_545));
	NAND2_X1_LVT multiplier_0i_32_500 (.A1(multiplier_0_n_32_33),.A2(multiplier_0_n_32_545),.ZN(multiplier_0_n_32_544));
	NAND2_X1_LVT multiplier_0i_32_48 (.A1(multiplier_0_op2_xp[2]),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_32_48));
	NAND2_X1_LVT multiplier_0i_32_64 (.A1(multiplier_0_op2_xp[3]),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_32_64));
	NOR2_X1_LVT multiplier_0i_32_473 (.A1(multiplier_0_n_32_48),.A2(multiplier_0_n_32_64),.ZN(multiplier_0_n_32_512));
	NAND2_X1_LVT multiplier_0i_32_32 (.A1(multiplier_0_op2_xp[1]),.A2(multiplier_0_op1[15]),.ZN(multiplier_0_n_32_32));
	NOR2_X1_LVT multiplier_0i_32_474 (.A1(multiplier_0_n_32_32),.A2(multiplier_0_n_32_64),.ZN(multiplier_0_n_32_513));
	NOR2_X1_LVT multiplier_0i_32_475 (.A1(multiplier_0_n_32_32),.A2(multiplier_0_n_32_48),.ZN(multiplier_0_n_32_514));
	OR3_X1_LVT multiplier_0i_32_472 (.A1(multiplier_0_n_32_512),.A2(multiplier_0_n_32_513),.A3(multiplier_0_n_32_514),.ZN(multiplier_0_n_32_511));
	NAND2_X1_LVT multiplier_0i_32_502 (.A1(multiplier_0_n_32_511),.A2(multiplier_0_n_32_545),.ZN(multiplier_0_n_32_546));
	NAND2_X1_LVT multiplier_0i_32_503 (.A1(multiplier_0_n_32_511),.A2(multiplier_0_n_32_33),.ZN(multiplier_0_n_32_547));
	NAND3_X1_LVT multiplier_0i_32_499 (.A1(multiplier_0_n_32_544),.A2(multiplier_0_n_32_546),.A3(multiplier_0_n_32_547),.ZN(multiplier_0_n_32_543));
	NAND2_X1_LVT multiplier_0i_32_96 (.A1(multiplier_0_op2_xp[5]),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_32_96));
	NAND2_X1_LVT multiplier_0i_32_112 (.A1(multiplier_0_op2_xp[6]),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_32_112));
	NOR2_X1_LVT multiplier_0i_32_466 (.A1(multiplier_0_n_32_96),.A2(multiplier_0_n_32_112),.ZN(multiplier_0_n_32_505));
	NAND2_X1_LVT multiplier_0i_32_80 (.A1(multiplier_0_op2_xp[4]),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_32_80));
	NOR2_X1_LVT multiplier_0i_32_467 (.A1(multiplier_0_n_32_80),.A2(multiplier_0_n_32_112),.ZN(multiplier_0_n_32_506));
	NOR2_X1_LVT multiplier_0i_32_468 (.A1(multiplier_0_n_32_80),.A2(multiplier_0_n_32_96),.ZN(multiplier_0_n_32_507));
	OR3_X1_LVT multiplier_0i_32_465 (.A1(multiplier_0_n_32_505),.A2(multiplier_0_n_32_506),.A3(multiplier_0_n_32_507),.ZN(multiplier_0_n_32_504));
	NAND2_X1_LVT multiplier_0i_32_128 (.A1(multiplier_0_op2_xp[7]),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_32_128));
	NAND2_X1_LVT multiplier_0i_32_144 (.A1(multiplier_0_op2_xp[8]),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_32_144));
	INV_X1_LVT multiplier_0i_32_461 (.A(multiplier_0_n_32_144),.ZN(multiplier_0_n_32_500));
	NAND2_X1_LVT multiplier_0i_32_460 (.A1(multiplier_0_n_32_128),.A2(multiplier_0_n_32_500),.ZN(multiplier_0_n_32_499));
	NAND2_X1_LVT multiplier_0i_32_16 (.A1(multiplier_0_op2_xp[0]),.A2(multiplier_0_op1_xp[0]),.ZN(multiplier_0_n_32_16));
	NOR2_X1_LVT multiplier_0i_32_451 (.A1(multiplier_0_n_32_31),.A2(multiplier_0_n_32_47),.ZN(multiplier_0_n_32_486));
	NOR2_X1_LVT multiplier_0i_32_452 (.A1(multiplier_0_n_32_15),.A2(multiplier_0_n_32_47),.ZN(multiplier_0_n_32_487));
	NOR2_X1_LVT multiplier_0i_32_453 (.A1(multiplier_0_n_32_15),.A2(multiplier_0_n_32_31),.ZN(multiplier_0_n_32_488));
	OR3_X1_LVT multiplier_0i_32_450 (.A1(multiplier_0_n_32_486),.A2(multiplier_0_n_32_487),.A3(multiplier_0_n_32_488),.ZN(multiplier_0_n_32_485));
	NOR2_X1_LVT multiplier_0i_32_444 (.A1(multiplier_0_n_32_79),.A2(multiplier_0_n_32_95),.ZN(multiplier_0_n_32_479));
	NOR2_X1_LVT multiplier_0i_32_445 (.A1(multiplier_0_n_32_63),.A2(multiplier_0_n_32_95),.ZN(multiplier_0_n_32_480));
	NOR2_X1_LVT multiplier_0i_32_446 (.A1(multiplier_0_n_32_63),.A2(multiplier_0_n_32_79),.ZN(multiplier_0_n_32_481));
	OR3_X1_LVT multiplier_0i_32_443 (.A1(multiplier_0_n_32_479),.A2(multiplier_0_n_32_480),.A3(multiplier_0_n_32_481),.ZN(multiplier_0_n_32_478));
	FA_X1_LVT multiplier_0i_32_476 (.A(multiplier_0_n_32_16),.B(multiplier_0_n_32_485),.CI(multiplier_0_n_32_478),.CO(multiplier_0_n_32_516),.S(multiplier_0_n_32_515));
	FA_X1_LVT multiplier_0i_32_504 (.A(multiplier_0_n_32_504),.B(multiplier_0_n_32_499),.CI(multiplier_0_n_32_516),.CO(multiplier_0_n_32_549),.S(multiplier_0_n_32_548));
	XNOR2_X1_LVT multiplier_0i_32_516 (.A(multiplier_0_n_32_98),.B(multiplier_0_n_32_82),.ZN(multiplier_0_n_32_564));
	XNOR2_X1_LVT multiplier_0i_32_517 (.A(multiplier_0_n_32_564),.B(multiplier_0_n_32_66),.ZN(multiplier_0_n_32_565));
	INV_X1_LVT multiplier_0i_32_518 (.A(multiplier_0_n_32_565),.ZN(multiplier_0_n_32_566));
	FA_X1_LVT multiplier_0i_32_524 (.A(multiplier_0_n_32_543),.B(multiplier_0_n_32_549),.CI(multiplier_0_n_32_566),.CO(multiplier_0_n_32_574),.S(multiplier_0_n_32_573));
	XNOR2_X1_LVT multiplier_0i_32_508 (.A(multiplier_0_n_32_146),.B(multiplier_0_n_32_130),.ZN(multiplier_0_n_32_556));
	XNOR2_X1_LVT multiplier_0i_32_509 (.A(multiplier_0_n_32_556),.B(multiplier_0_n_32_114),.ZN(multiplier_0_n_32_557));
	XNOR2_X1_LVT multiplier_0i_32_496 (.A(multiplier_0_n_32_49),.B(multiplier_0_n_32_33),.ZN(multiplier_0_n_32_540));
	XNOR2_X1_LVT multiplier_0i_32_497 (.A(multiplier_0_n_32_540),.B(multiplier_0_n_32_511),.ZN(multiplier_0_n_32_541));
	INV_X1_LVT multiplier_0i_32_498 (.A(multiplier_0_n_32_541),.ZN(multiplier_0_n_32_542));
	XNOR2_X1_LVT multiplier_0i_32_489 (.A(multiplier_0_n_32_97),.B(multiplier_0_n_32_81),.ZN(multiplier_0_n_32_533));
	XNOR2_X1_LVT multiplier_0i_32_490 (.A(multiplier_0_n_32_533),.B(multiplier_0_n_32_65),.ZN(multiplier_0_n_32_534));
	INV_X1_LVT multiplier_0i_32_491 (.A(multiplier_0_n_32_534),.ZN(multiplier_0_n_32_535));
	XNOR2_X1_LVT multiplier_0i_32_481 (.A(multiplier_0_n_32_145),.B(multiplier_0_n_32_129),.ZN(multiplier_0_n_32_525));
	XNOR2_X1_LVT multiplier_0i_32_482 (.A(multiplier_0_n_32_525),.B(multiplier_0_n_32_113),.ZN(multiplier_0_n_32_526));
	FA_X1_LVT multiplier_0i_32_505 (.A(multiplier_0_n_32_542),.B(multiplier_0_n_32_535),.CI(multiplier_0_n_32_526),.CO(multiplier_0_n_32_551),.S(multiplier_0_n_32_550));
	FA_X1_LVT multiplier_0i_32_525 (.A(multiplier_0_n_32_557),.B(multiplier_0_n_32_571),.CI(multiplier_0_n_32_551),.CO(multiplier_0_n_32_576),.S(multiplier_0_n_32_575));
	FA_X1_LVT multiplier_0i_32_545 (.A(multiplier_0_n_32_574),.B(multiplier_0_n_32_576),.CI(multiplier_0_n_32_597),.CO(multiplier_0_n_32_600),.S(multiplier_0_n_32_599));
	INV_X1_LVT multiplier_0i_32_436 (.A(multiplier_0_n_32_127),.ZN(multiplier_0_n_32_471));
	NAND2_X1_LVT multiplier_0i_32_435 (.A1(multiplier_0_n_32_143),.A2(multiplier_0_n_32_471),.ZN(multiplier_0_n_32_470));
	INV_X1_LVT multiplier_0i_32_438 (.A(multiplier_0_n_32_111),.ZN(multiplier_0_n_32_473));
	NAND2_X1_LVT multiplier_0i_32_437 (.A1(multiplier_0_n_32_143),.A2(multiplier_0_n_32_473),.ZN(multiplier_0_n_32_472));
	OR2_X1_LVT multiplier_0i_32_439 (.A1(multiplier_0_n_32_111),.A2(multiplier_0_n_32_127),.ZN(multiplier_0_n_32_474));
	NAND3_X1_LVT multiplier_0i_32_434 (.A1(multiplier_0_n_32_470),.A2(multiplier_0_n_32_472),.A3(multiplier_0_n_32_474),.ZN(multiplier_0_n_32_469));
	XNOR2_X1_LVT multiplier_0i_32_469 (.A(multiplier_0_n_32_64),.B(multiplier_0_n_32_48),.ZN(multiplier_0_n_32_508));
	XNOR2_X1_LVT multiplier_0i_32_470 (.A(multiplier_0_n_32_508),.B(multiplier_0_n_32_32),.ZN(multiplier_0_n_32_509));
	INV_X1_LVT multiplier_0i_32_471 (.A(multiplier_0_n_32_509),.ZN(multiplier_0_n_32_510));
	FA_X1_LVT multiplier_0i_32_477 (.A(multiplier_0_n_32_469),.B(multiplier_0_n_32_490),.CI(multiplier_0_n_32_510),.CO(multiplier_0_n_32_518),.S(multiplier_0_n_32_517));
	XNOR2_X1_LVT multiplier_0i_32_462 (.A(multiplier_0_n_32_112),.B(multiplier_0_n_32_96),.ZN(multiplier_0_n_32_501));
	XNOR2_X1_LVT multiplier_0i_32_463 (.A(multiplier_0_n_32_501),.B(multiplier_0_n_32_80),.ZN(multiplier_0_n_32_502));
	INV_X1_LVT multiplier_0i_32_464 (.A(multiplier_0_n_32_502),.ZN(multiplier_0_n_32_503));
	XNOR2_X1_LVT multiplier_0i_32_458 (.A(multiplier_0_n_32_144),.B(multiplier_0_n_32_128),.ZN(multiplier_0_n_32_497));
	INV_X1_LVT multiplier_0i_32_459 (.A(multiplier_0_n_32_497),.ZN(multiplier_0_n_32_498));
	FA_X1_LVT multiplier_0i_32_478 (.A(multiplier_0_n_32_503),.B(multiplier_0_n_32_498),.CI(multiplier_0_n_32_515),.CO(multiplier_0_n_32_520),.S(multiplier_0_n_32_519));
	FA_X1_LVT multiplier_0i_32_506 (.A(multiplier_0_n_32_548),.B(multiplier_0_n_32_518),.CI(multiplier_0_n_32_520),.CO(multiplier_0_n_32_553),.S(multiplier_0_n_32_552));
	FA_X1_LVT multiplier_0i_32_526 (.A(multiplier_0_n_32_573),.B(multiplier_0_n_32_553),.CI(multiplier_0_n_32_575),.CO(multiplier_0_n_32_578),.S(multiplier_0_n_32_577));
	FA_X1_LVT multiplier_0i_32_479 (.A(multiplier_0_n_32_492),.B(multiplier_0_n_32_517),.CI(multiplier_0_n_32_494),.CO(multiplier_0_n_32_522),.S(multiplier_0_n_32_521));
	FA_X1_LVT multiplier_0i_32_507 (.A(multiplier_0_n_32_522),.B(multiplier_0_n_32_550),.CI(multiplier_0_n_32_552),.CO(multiplier_0_n_32_555),.S(multiplier_0_n_32_554));
	HA_X1_LVT multiplier_0i_32_480 (.A(multiplier_0_n_32_519),.B(multiplier_0_n_32_521),.CO(multiplier_0_n_32_524),.S(multiplier_0_n_32_523));
	FA_X1_LVT multiplier_0i_32_610 (.A(multiplier_0_n_32_496),.B(multiplier_0_n_32_523),.CI(multiplier_0_n_32_666),.CO(multiplier_0_n_32_667),.S(multiplier_0_n_58));
	FA_X1_LVT multiplier_0i_32_611 (.A(multiplier_0_n_32_524),.B(multiplier_0_n_32_554),.CI(multiplier_0_n_32_667),.CO(multiplier_0_n_32_668),.S(multiplier_0_n_59));
	FA_X1_LVT multiplier_0i_32_612 (.A(multiplier_0_n_32_555),.B(multiplier_0_n_32_577),.CI(multiplier_0_n_32_668),.CO(multiplier_0_n_32_669),.S(multiplier_0_n_60));
	FA_X1_LVT multiplier_0i_32_613 (.A(multiplier_0_n_32_599),.B(multiplier_0_n_32_578),.CI(multiplier_0_n_32_669),.CO(multiplier_0_n_32_670),.S(multiplier_0_n_61));
	FA_X1_LVT multiplier_0i_32_614 (.A(multiplier_0_n_32_600),.B(multiplier_0_n_32_619),.CI(multiplier_0_n_32_670),.CO(multiplier_0_n_32_671),.S(multiplier_0_n_62));
	FA_X1_LVT multiplier_0i_32_615 (.A(multiplier_0_n_32_620),.B(multiplier_0_n_32_631),.CI(multiplier_0_n_32_671),.CO(multiplier_0_n_32_672),.S(multiplier_0_n_63));
	FA_X1_LVT multiplier_0i_32_616 (.A(multiplier_0_n_32_632),.B(multiplier_0_n_32_641),.CI(multiplier_0_n_32_672),.CO(multiplier_0_n_32_673),.S(multiplier_0_n_64));
	XNOR2_X1_LVT multiplier_0i_32_618 (.A(multiplier_0_n_32_674),.B(multiplier_0_n_32_673),.ZN(multiplier_0_n_65));
	AND2_X1_LVT multiplier_0i_33_0 (.A1(multiplier_0_sign_sel),.A2(multiplier_0_n_65),.ZN(multiplier_0_n_66));
	NAND2_X1_LVT multiplier_0i_34_49 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_66),.ZN(multiplier_0_n_34_25));
	INV_X1_LVT multiplier_0i_34_47 (.A(multiplier_0_n_65),.ZN(multiplier_0_n_34_24));
	OAI21_X1_LVT multiplier_0i_34_57 (.A(multiplier_0_n_34_25),.B1(multiplier_0_n_34_8),.B2(multiplier_0_n_34_24),.ZN(multiplier_0_product_xp[0]));
	NOR3_X1_LVT multiplier_0i_3_9 (.A1(multiplier_0_n_3_2),.A2(multiplier_0_n_3_1),.A3(per_addr[0]),.ZN(multiplier_0_n_7));
	AND2_X1_LVT multiplier_0i_7_6 (.A1(multiplier_0_reg_write),.A2(multiplier_0_n_7),.ZN(multiplier_0_reshi_wr));
	NOR2_X1_LVT multiplier_0i_41_0 (.A1(multiplier_0_result_clr),.A2(multiplier_0_reshi_wr),.ZN(multiplier_0_n_41_0));
	AOI22_X1_LVT multiplier_0i_41_31 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[15]),.B1(multiplier_0_reshi_wr),.B2(multiplier_0_per_din_msk[15]),.ZN(multiplier_0_n_41_16));
	INV_X1_LVT multiplier_0i_41_32 (.A(multiplier_0_n_41_16),.ZN(multiplier_0_n_86));
	INV_X1_LVT multiplier_0i_42_1 (.A(multiplier_0_n_69),.ZN(multiplier_0_n_42_1));
	INV_X1_LVT multiplier_0i_42_0 (.A(multiplier_0_reshi_wr),.ZN(multiplier_0_n_42_0));
	NAND2_X1_LVT multiplier_0i_42_2 (.A1(multiplier_0_n_42_1),.A2(multiplier_0_n_42_0),.ZN(multiplier_0_n_87));
	CLKGATETST_X1_LVT multiplier_0clk_gate_reshi_reg (.CK(mclk),.E(multiplier_0_n_87),.SE(1'b0),.GCK(multiplier_0_n_70));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b15___05F05d (.D(multiplier_0_n_86),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[15]),.QN());
	INV_X1_LVT multiplier_0i_34_45 (.A(multiplier_0_n_64),.ZN(multiplier_0_n_34_23));
	OAI21_X1_LVT multiplier_0i_34_56 (.A(multiplier_0_n_34_25),.B1(multiplier_0_n_34_8),.B2(multiplier_0_n_34_23),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_29 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[14]),.B1(multiplier_0_reshi_wr),.B2(multiplier_0_per_din_msk[14]),.ZN(multiplier_0_n_41_15));
	INV_X1_LVT multiplier_0i_41_30 (.A(multiplier_0_n_41_15),.ZN(multiplier_0_n_85));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b14___05F05d (.D(multiplier_0_n_85),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[14]),.QN());
	INV_X1_LVT multiplier_0i_34_43 (.A(multiplier_0_n_63),.ZN(multiplier_0_n_34_22));
	OAI21_X1_LVT multiplier_0i_34_55 (.A(multiplier_0_n_34_25),.B1(multiplier_0_n_34_8),.B2(multiplier_0_n_34_22),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_27 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[13]),.B1(multiplier_0_reshi_wr),.B2(multiplier_0_per_din_msk[13]),.ZN(multiplier_0_n_41_14));
	INV_X1_LVT multiplier_0i_41_28 (.A(multiplier_0_n_41_14),.ZN(multiplier_0_n_84));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b13___05F05d (.D(multiplier_0_n_84),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[13]),.QN());
	INV_X1_LVT multiplier_0i_34_41 (.A(multiplier_0_n_62),.ZN(multiplier_0_n_34_21));
	OAI21_X1_LVT multiplier_0i_34_54 (.A(multiplier_0_n_34_25),.B1(multiplier_0_n_34_8),.B2(multiplier_0_n_34_21),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_25 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[12]),.B1(multiplier_0_reshi_wr),.B2(multiplier_0_per_din_msk[12]),.ZN(multiplier_0_n_41_13));
	INV_X1_LVT multiplier_0i_41_26 (.A(multiplier_0_n_41_13),.ZN(multiplier_0_n_83));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b12___05F05d (.D(multiplier_0_n_83),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[12]),.QN());
	INV_X1_LVT multiplier_0i_34_39 (.A(multiplier_0_n_61),.ZN(multiplier_0_n_34_20));
	OAI21_X1_LVT multiplier_0i_34_53 (.A(multiplier_0_n_34_25),.B1(multiplier_0_n_34_8),.B2(multiplier_0_n_34_20),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_23 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[11]),.B1(multiplier_0_reshi_wr),.B2(multiplier_0_per_din_msk[11]),.ZN(multiplier_0_n_41_12));
	INV_X1_LVT multiplier_0i_41_24 (.A(multiplier_0_n_41_12),.ZN(multiplier_0_n_82));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b11___05F05d (.D(multiplier_0_n_82),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[11]),.QN());
	INV_X1_LVT multiplier_0i_34_37 (.A(multiplier_0_n_60),.ZN(multiplier_0_n_34_19));
	OAI21_X1_LVT multiplier_0i_34_52 (.A(multiplier_0_n_34_25),.B1(multiplier_0_n_34_8),.B2(multiplier_0_n_34_19),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_21 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[10]),.B1(multiplier_0_reshi_wr),.B2(multiplier_0_per_din_msk[10]),.ZN(multiplier_0_n_41_11));
	INV_X1_LVT multiplier_0i_41_22 (.A(multiplier_0_n_41_11),.ZN(multiplier_0_n_81));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b10___05F05d (.D(multiplier_0_n_81),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[10]),.QN());
	INV_X1_LVT multiplier_0i_34_35 (.A(multiplier_0_n_59),.ZN(multiplier_0_n_34_18));
	OAI21_X1_LVT multiplier_0i_34_51 (.A(multiplier_0_n_34_25),.B1(multiplier_0_n_34_8),.B2(multiplier_0_n_34_18),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_19 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[9]),.B1(multiplier_0_reshi_wr),.B2(multiplier_0_per_din_msk[9]),.ZN(multiplier_0_n_41_10));
	INV_X1_LVT multiplier_0i_41_20 (.A(multiplier_0_n_41_10),.ZN(multiplier_0_n_80));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b9___05F05d (.D(multiplier_0_n_80),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[9]),.QN());
	INV_X1_LVT multiplier_0i_34_33 (.A(multiplier_0_n_58),.ZN(multiplier_0_n_34_17));
	OAI21_X1_LVT multiplier_0i_34_50 (.A(multiplier_0_n_34_25),.B1(multiplier_0_n_34_8),.B2(multiplier_0_n_34_17),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_17 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[8]),.B1(multiplier_0_reshi_wr),.B2(multiplier_0_per_din_msk[8]),.ZN(multiplier_0_n_41_9));
	INV_X1_LVT multiplier_0i_41_18 (.A(multiplier_0_n_41_9),.ZN(multiplier_0_n_79));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b8___05F05d (.D(multiplier_0_n_79),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[8]),.QN());
	OAI22_X1_LVT multiplier_0i_34_48 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_16),.B1(multiplier_0_n_34_24),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_15 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[7]),.B1(multiplier_0_reshi_wr),.B2(per_din[7]),.ZN(multiplier_0_n_41_8));
	INV_X1_LVT multiplier_0i_41_16 (.A(multiplier_0_n_41_8),.ZN(multiplier_0_n_78));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b7___05F05d (.D(multiplier_0_n_78),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[7]),.QN());
	OAI22_X1_LVT multiplier_0i_34_46 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_15),.B1(multiplier_0_n_34_23),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_13 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[6]),.B1(multiplier_0_reshi_wr),.B2(per_din[6]),.ZN(multiplier_0_n_41_7));
	INV_X1_LVT multiplier_0i_41_14 (.A(multiplier_0_n_41_7),.ZN(multiplier_0_n_77));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b6___05F05d (.D(multiplier_0_n_77),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[6]),.QN());
	OAI22_X1_LVT multiplier_0i_34_44 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_14),.B1(multiplier_0_n_34_22),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_11 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[5]),.B1(multiplier_0_reshi_wr),.B2(per_din[5]),.ZN(multiplier_0_n_41_6));
	INV_X1_LVT multiplier_0i_41_12 (.A(multiplier_0_n_41_6),.ZN(multiplier_0_n_76));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b5___05F05d (.D(multiplier_0_n_76),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[5]),.QN());
	OAI22_X1_LVT multiplier_0i_34_42 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_13),.B1(multiplier_0_n_34_21),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_9 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[4]),.B1(multiplier_0_reshi_wr),.B2(per_din[4]),.ZN(multiplier_0_n_41_5));
	INV_X1_LVT multiplier_0i_41_10 (.A(multiplier_0_n_41_5),.ZN(multiplier_0_n_75));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b4___05F05d (.D(multiplier_0_n_75),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[4]),.QN());
	OAI22_X1_LVT multiplier_0i_34_40 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_12),.B1(multiplier_0_n_34_20),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_7 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[3]),.B1(multiplier_0_reshi_wr),.B2(per_din[3]),.ZN(multiplier_0_n_41_4));
	INV_X1_LVT multiplier_0i_41_8 (.A(multiplier_0_n_41_4),.ZN(multiplier_0_n_74));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b3___05F05d (.D(multiplier_0_n_74),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[3]),.QN());
	OAI22_X1_LVT multiplier_0i_34_38 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_11),.B1(multiplier_0_n_34_19),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_5 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[2]),.B1(multiplier_0_reshi_wr),.B2(per_din[2]),.ZN(multiplier_0_n_41_3));
	INV_X1_LVT multiplier_0i_41_6 (.A(multiplier_0_n_41_3),.ZN(multiplier_0_n_73));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b2___05F05d (.D(multiplier_0_n_73),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[2]),.QN());
	OAI22_X1_LVT multiplier_0i_34_36 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_10),.B1(multiplier_0_n_34_18),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_3 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[1]),.B1(multiplier_0_reshi_wr),.B2(per_din[1]),.ZN(multiplier_0_n_41_2));
	INV_X1_LVT multiplier_0i_41_4 (.A(multiplier_0_n_41_2),.ZN(multiplier_0_n_72));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b1___05F05d (.D(multiplier_0_n_72),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[1]),.QN());
	OAI22_X1_LVT multiplier_0i_34_34 (.A1(multiplier_0_n_34_8),.A2(multiplier_0_n_34_9),.B1(multiplier_0_n_34_17),.B2(multiplier_0_cycle[0]),.ZN(multiplier_0_product_xp[0]));
	AOI22_X1_LVT multiplier_0i_41_1 (.A1(multiplier_0_n_41_0),.A2(multiplier_0_reshi_nxt[0]),.B1(per_din[0]),.B2(multiplier_0_reshi_wr),.ZN(multiplier_0_n_41_1));
	INV_X1_LVT multiplier_0i_41_2 (.A(multiplier_0_n_41_1),.ZN(multiplier_0_n_71));
	DFFR_X1_LVT multiplier_0reshi_reg___05F05b0___05F05d (.D(multiplier_0_n_71),.RN(multiplier_0_n_38),.CK(multiplier_0_n_70),.Q(multiplier_0_reshi[0]),.QN());
	FA_X1_LVT multiplier_0i_48_16 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[0]),.CI(multiplier_0_n_48_15),.CO(multiplier_0_n_48_16),.S(multiplier_0_reshi_nxt[0]));
	FA_X1_LVT multiplier_0i_48_17 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[1]),.CI(multiplier_0_n_48_16),.CO(multiplier_0_n_48_17),.S(multiplier_0_reshi_nxt[1]));
	FA_X1_LVT multiplier_0i_48_18 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[2]),.CI(multiplier_0_n_48_17),.CO(multiplier_0_n_48_18),.S(multiplier_0_reshi_nxt[2]));
	FA_X1_LVT multiplier_0i_48_19 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[3]),.CI(multiplier_0_n_48_18),.CO(multiplier_0_n_48_19),.S(multiplier_0_reshi_nxt[3]));
	FA_X1_LVT multiplier_0i_48_20 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[4]),.CI(multiplier_0_n_48_19),.CO(multiplier_0_n_48_20),.S(multiplier_0_reshi_nxt[4]));
	FA_X1_LVT multiplier_0i_48_21 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[5]),.CI(multiplier_0_n_48_20),.CO(multiplier_0_n_48_21),.S(multiplier_0_reshi_nxt[5]));
	FA_X1_LVT multiplier_0i_48_22 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[6]),.CI(multiplier_0_n_48_21),.CO(multiplier_0_n_48_22),.S(multiplier_0_reshi_nxt[6]));
	FA_X1_LVT multiplier_0i_48_23 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[7]),.CI(multiplier_0_n_48_22),.CO(multiplier_0_n_48_23),.S(multiplier_0_reshi_nxt[7]));
	FA_X1_LVT multiplier_0i_48_24 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[8]),.CI(multiplier_0_n_48_23),.CO(multiplier_0_n_48_24),.S(multiplier_0_reshi_nxt[8]));
	FA_X1_LVT multiplier_0i_48_25 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[9]),.CI(multiplier_0_n_48_24),.CO(multiplier_0_n_48_25),.S(multiplier_0_reshi_nxt[9]));
	FA_X1_LVT multiplier_0i_48_26 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[10]),.CI(multiplier_0_n_48_25),.CO(multiplier_0_n_48_26),.S(multiplier_0_reshi_nxt[10]));
	FA_X1_LVT multiplier_0i_48_27 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[11]),.CI(multiplier_0_n_48_26),.CO(multiplier_0_n_48_27),.S(multiplier_0_reshi_nxt[11]));
	FA_X1_LVT multiplier_0i_48_28 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[12]),.CI(multiplier_0_n_48_27),.CO(multiplier_0_n_48_28),.S(multiplier_0_reshi_nxt[12]));
	FA_X1_LVT multiplier_0i_48_29 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[13]),.CI(multiplier_0_n_48_28),.CO(multiplier_0_n_48_29),.S(multiplier_0_reshi_nxt[13]));
	FA_X1_LVT multiplier_0i_48_30 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[14]),.CI(multiplier_0_n_48_29),.CO(multiplier_0_n_48_30),.S(multiplier_0_reshi_nxt[14]));
	FA_X1_LVT multiplier_0i_48_31 (.A(multiplier_0_product_xp[0]),.B(multiplier_0_reshi[15]),.CI(multiplier_0_n_48_30),.CO(multiplier_0_n_138),.S(multiplier_0_reshi_nxt[15]));
	NAND2_X1_LVT multiplier_0i_50_0 (.A1(multiplier_0_reshi_nxt[15]),.A2(multiplier_0_sign_sel),.ZN(multiplier_0_n_50_0));
	INV_X1_LVT multiplier_0i_50_3 (.A(multiplier_0_n_50_0),.ZN(multiplier_0_sumext_s_nxt[1]));
	AND2_X1_LVT multiplier_0i_52_2 (.A1(multiplier_0_n_52_0),.A2(multiplier_0_sumext_s_nxt[1]),.ZN(multiplier_0_n_142));
	INV_X1_LVT multiplier_0i_53_1 (.A(multiplier_0_result_wr),.ZN(multiplier_0_n_53_1));
	INV_X1_LVT multiplier_0i_53_0 (.A(multiplier_0_op2_wr),.ZN(multiplier_0_n_53_0));
	NAND2_X1_LVT multiplier_0i_53_2 (.A1(multiplier_0_n_53_1),.A2(multiplier_0_n_53_0),.ZN(multiplier_0_n_143));
	CLKGATETST_X1_LVT multiplier_0clk_gate_sumext_s_reg (.CK(mclk),.E(multiplier_0_n_143),.SE(1'b0),.GCK(multiplier_0_n_140));
	DFFR_X1_LVT multiplier_0sumext_s_reg___05F05b1___05F05d (.D(multiplier_0_n_142),.RN(multiplier_0_n_38),.CK(multiplier_0_n_140),.Q(multiplier_0_sumext_s[1]),.QN());
	AOI22_X1_LVT multiplier_0i_57_1 (.A1(multiplier_0_n_57_0),.A2(multiplier_0_sumext_s[1]),.B1(multiplier_0_sumext_s_nxt[1]),.B2(multiplier_0_cycle[1]),.ZN(multiplier_0_n_57_1));
	INV_X1_LVT multiplier_0i_57_2 (.A(multiplier_0_n_57_1),.ZN(multiplier_0_n_148));
	NOR3_X1_LVT multiplier_0i_3_10 (.A1(multiplier_0_n_3_0),.A2(multiplier_0_n_3_1),.A3(multiplier_0_n_3_2),.ZN(multiplier_0_n_8));
	AND2_X1_LVT multiplier_0i_4_7 (.A1(multiplier_0_reg_read),.A2(multiplier_0_n_8),.ZN(multiplier_0_reg_rd15));
	AND2_X1_LVT multiplier_0i_58_0 (.A1(multiplier_0_n_148),.A2(multiplier_0_reg_rd15),.ZN(multiplier_0_n_149));
	AND2_X1_LVT multiplier_0i_4_4 (.A1(multiplier_0_reg_read),.A2(multiplier_0_n_5),.ZN(multiplier_0_n_12));
	AND2_X1_LVT multiplier_0i_20_0 (.A1(multiplier_0_op2_reg[15]),.A2(multiplier_0_n_12),.ZN(multiplier_0_n_37));
	NOR4_X1_LVT multiplier_0i_60_96 (.A1(multiplier_0_n_60_79),.A2(multiplier_0_n_60_80),.A3(multiplier_0_n_149),.A4(multiplier_0_n_37),.ZN(multiplier_0_n_60_81));
	AOI22_X1_LVT multiplier_0i_60_97 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[15]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[15]),.ZN(multiplier_0_n_60_82));
	AND2_X1_LVT multiplier_0i_4_6 (.A1(multiplier_0_reg_read),.A2(multiplier_0_n_7),.ZN(multiplier_0_n_14));
	INV_X1_LVT multiplier_0i_60_7 (.A(multiplier_0_n_14),.ZN(multiplier_0_n_60_7));
	OAI21_X1_LVT multiplier_0i_60_98 (.A(multiplier_0_n_60_81),.B1(multiplier_0_n_60_82),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[15]));
	AOI22_X1_LVT multiplier_0i_60_87 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_90),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_136),.ZN(multiplier_0_n_60_73));
	NOR2_X1_LVT multiplier_0i_60_88 (.A1(multiplier_0_n_60_73),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_74));
	AND2_X1_LVT multiplier_0i_60_89 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[14]),.ZN(multiplier_0_n_60_75));
	AND2_X1_LVT multiplier_0i_19_0 (.A1(multiplier_0_op2_reg[14]),.A2(multiplier_0_n_12),.ZN(multiplier_0_n_36));
	NOR4_X1_LVT multiplier_0i_60_90 (.A1(multiplier_0_n_60_74),.A2(multiplier_0_n_60_75),.A3(multiplier_0_n_149),.A4(multiplier_0_n_36),.ZN(multiplier_0_n_60_76));
	AOI22_X1_LVT multiplier_0i_60_91 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[14]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[14]),.ZN(multiplier_0_n_60_77));
	OAI21_X1_LVT multiplier_0i_60_92 (.A(multiplier_0_n_60_76),.B1(multiplier_0_n_60_77),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[14]));
	AOI22_X1_LVT multiplier_0i_60_81 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_91),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_135),.ZN(multiplier_0_n_60_68));
	NOR2_X1_LVT multiplier_0i_60_82 (.A1(multiplier_0_n_60_68),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_69));
	AND2_X1_LVT multiplier_0i_60_83 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[13]),.ZN(multiplier_0_n_60_70));
	AND2_X1_LVT multiplier_0i_18_0 (.A1(multiplier_0_op2_reg[13]),.A2(multiplier_0_n_12),.ZN(multiplier_0_n_35));
	NOR4_X1_LVT multiplier_0i_60_84 (.A1(multiplier_0_n_60_69),.A2(multiplier_0_n_60_70),.A3(multiplier_0_n_149),.A4(multiplier_0_n_35),.ZN(multiplier_0_n_60_71));
	AOI22_X1_LVT multiplier_0i_60_85 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[13]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[13]),.ZN(multiplier_0_n_60_72));
	OAI21_X1_LVT multiplier_0i_60_86 (.A(multiplier_0_n_60_71),.B1(multiplier_0_n_60_72),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[13]));
	AOI22_X1_LVT multiplier_0i_60_75 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_92),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_134),.ZN(multiplier_0_n_60_63));
	NOR2_X1_LVT multiplier_0i_60_76 (.A1(multiplier_0_n_60_63),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_64));
	AND2_X1_LVT multiplier_0i_60_77 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[12]),.ZN(multiplier_0_n_60_65));
	AND2_X1_LVT multiplier_0i_17_0 (.A1(multiplier_0_op2_reg[12]),.A2(multiplier_0_n_12),.ZN(multiplier_0_n_34));
	NOR4_X1_LVT multiplier_0i_60_78 (.A1(multiplier_0_n_60_64),.A2(multiplier_0_n_60_65),.A3(multiplier_0_n_149),.A4(multiplier_0_n_34),.ZN(multiplier_0_n_60_66));
	AOI22_X1_LVT multiplier_0i_60_79 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[12]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[12]),.ZN(multiplier_0_n_60_67));
	OAI21_X1_LVT multiplier_0i_60_80 (.A(multiplier_0_n_60_66),.B1(multiplier_0_n_60_67),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[12]));
	AOI22_X1_LVT multiplier_0i_60_69 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_93),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_133),.ZN(multiplier_0_n_60_58));
	NOR2_X1_LVT multiplier_0i_60_70 (.A1(multiplier_0_n_60_58),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_59));
	AND2_X1_LVT multiplier_0i_60_71 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[11]),.ZN(multiplier_0_n_60_60));
	AND2_X1_LVT multiplier_0i_16_0 (.A1(multiplier_0_op2_reg[11]),.A2(multiplier_0_n_12),.ZN(multiplier_0_n_33));
	NOR4_X1_LVT multiplier_0i_60_72 (.A1(multiplier_0_n_60_59),.A2(multiplier_0_n_60_60),.A3(multiplier_0_n_149),.A4(multiplier_0_n_33),.ZN(multiplier_0_n_60_61));
	AOI22_X1_LVT multiplier_0i_60_73 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[11]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[11]),.ZN(multiplier_0_n_60_62));
	OAI21_X1_LVT multiplier_0i_60_74 (.A(multiplier_0_n_60_61),.B1(multiplier_0_n_60_62),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[11]));
	AOI22_X1_LVT multiplier_0i_60_63 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_94),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_132),.ZN(multiplier_0_n_60_53));
	NOR2_X1_LVT multiplier_0i_60_64 (.A1(multiplier_0_n_60_53),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_54));
	AND2_X1_LVT multiplier_0i_60_65 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[10]),.ZN(multiplier_0_n_60_55));
	AND2_X1_LVT multiplier_0i_15_0 (.A1(multiplier_0_op2_reg[10]),.A2(multiplier_0_n_12),.ZN(multiplier_0_n_32));
	NOR4_X1_LVT multiplier_0i_60_66 (.A1(multiplier_0_n_60_54),.A2(multiplier_0_n_60_55),.A3(multiplier_0_n_149),.A4(multiplier_0_n_32),.ZN(multiplier_0_n_60_56));
	AOI22_X1_LVT multiplier_0i_60_67 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[10]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[10]),.ZN(multiplier_0_n_60_57));
	OAI21_X1_LVT multiplier_0i_60_68 (.A(multiplier_0_n_60_56),.B1(multiplier_0_n_60_57),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[10]));
	AOI22_X1_LVT multiplier_0i_60_57 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_95),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_131),.ZN(multiplier_0_n_60_48));
	NOR2_X1_LVT multiplier_0i_60_58 (.A1(multiplier_0_n_60_48),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_49));
	AND2_X1_LVT multiplier_0i_60_59 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[9]),.ZN(multiplier_0_n_60_50));
	AND2_X1_LVT multiplier_0i_14_0 (.A1(multiplier_0_op2_reg[9]),.A2(multiplier_0_n_12),.ZN(multiplier_0_n_31));
	NOR4_X1_LVT multiplier_0i_60_60 (.A1(multiplier_0_n_60_49),.A2(multiplier_0_n_60_50),.A3(multiplier_0_n_149),.A4(multiplier_0_n_31),.ZN(multiplier_0_n_60_51));
	AOI22_X1_LVT multiplier_0i_60_61 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[9]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[9]),.ZN(multiplier_0_n_60_52));
	OAI21_X1_LVT multiplier_0i_60_62 (.A(multiplier_0_n_60_51),.B1(multiplier_0_n_60_52),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[9]));
	AOI22_X1_LVT multiplier_0i_60_51 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_96),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_130),.ZN(multiplier_0_n_60_43));
	NOR2_X1_LVT multiplier_0i_60_52 (.A1(multiplier_0_n_60_43),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_44));
	AND2_X1_LVT multiplier_0i_60_53 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[8]),.ZN(multiplier_0_n_60_45));
	AND2_X1_LVT multiplier_0i_13_0 (.A1(multiplier_0_op2_reg[8]),.A2(multiplier_0_n_12),.ZN(multiplier_0_n_30));
	NOR4_X1_LVT multiplier_0i_60_54 (.A1(multiplier_0_n_60_44),.A2(multiplier_0_n_60_45),.A3(multiplier_0_n_149),.A4(multiplier_0_n_30),.ZN(multiplier_0_n_60_46));
	AOI22_X1_LVT multiplier_0i_60_55 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[8]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[8]),.ZN(multiplier_0_n_60_47));
	OAI21_X1_LVT multiplier_0i_60_56 (.A(multiplier_0_n_60_46),.B1(multiplier_0_n_60_47),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[8]));
	AOI22_X1_LVT multiplier_0i_60_45 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_97),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_129),.ZN(multiplier_0_n_60_38));
	NOR2_X1_LVT multiplier_0i_60_46 (.A1(multiplier_0_n_60_38),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_39));
	AND2_X1_LVT multiplier_0i_60_47 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[7]),.ZN(multiplier_0_n_60_40));
	AND2_X1_LVT multiplier_0i_12_7 (.A1(multiplier_0_n_12),.A2(multiplier_0_op2_reg[7]),.ZN(multiplier_0_n_29));
	NOR4_X1_LVT multiplier_0i_60_48 (.A1(multiplier_0_n_60_39),.A2(multiplier_0_n_60_40),.A3(multiplier_0_n_149),.A4(multiplier_0_n_29),.ZN(multiplier_0_n_60_41));
	AOI22_X1_LVT multiplier_0i_60_49 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[7]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[7]),.ZN(multiplier_0_n_60_42));
	OAI21_X1_LVT multiplier_0i_60_50 (.A(multiplier_0_n_60_41),.B1(multiplier_0_n_60_42),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[7]));
	AOI22_X1_LVT multiplier_0i_60_39 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_98),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_128),.ZN(multiplier_0_n_60_33));
	NOR2_X1_LVT multiplier_0i_60_40 (.A1(multiplier_0_n_60_33),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_34));
	AND2_X1_LVT multiplier_0i_60_41 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[6]),.ZN(multiplier_0_n_60_35));
	AND2_X1_LVT multiplier_0i_12_6 (.A1(multiplier_0_n_12),.A2(multiplier_0_op2_reg[6]),.ZN(multiplier_0_n_28));
	NOR4_X1_LVT multiplier_0i_60_42 (.A1(multiplier_0_n_60_34),.A2(multiplier_0_n_60_35),.A3(multiplier_0_n_149),.A4(multiplier_0_n_28),.ZN(multiplier_0_n_60_36));
	AOI22_X1_LVT multiplier_0i_60_43 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[6]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[6]),.ZN(multiplier_0_n_60_37));
	OAI21_X1_LVT multiplier_0i_60_44 (.A(multiplier_0_n_60_36),.B1(multiplier_0_n_60_37),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[6]));
	AOI22_X1_LVT multiplier_0i_60_33 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_99),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_127),.ZN(multiplier_0_n_60_28));
	NOR2_X1_LVT multiplier_0i_60_34 (.A1(multiplier_0_n_60_28),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_29));
	AND2_X1_LVT multiplier_0i_60_35 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[5]),.ZN(multiplier_0_n_60_30));
	AND2_X1_LVT multiplier_0i_12_5 (.A1(multiplier_0_n_12),.A2(multiplier_0_op2_reg[5]),.ZN(multiplier_0_n_27));
	NOR4_X1_LVT multiplier_0i_60_36 (.A1(multiplier_0_n_60_29),.A2(multiplier_0_n_60_30),.A3(multiplier_0_n_149),.A4(multiplier_0_n_27),.ZN(multiplier_0_n_60_31));
	AOI22_X1_LVT multiplier_0i_60_37 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[5]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[5]),.ZN(multiplier_0_n_60_32));
	OAI21_X1_LVT multiplier_0i_60_38 (.A(multiplier_0_n_60_31),.B1(multiplier_0_n_60_32),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[5]));
	AOI22_X1_LVT multiplier_0i_60_27 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_100),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_126),.ZN(multiplier_0_n_60_23));
	NOR2_X1_LVT multiplier_0i_60_28 (.A1(multiplier_0_n_60_23),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_24));
	AND2_X1_LVT multiplier_0i_60_29 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[4]),.ZN(multiplier_0_n_60_25));
	AND2_X1_LVT multiplier_0i_12_4 (.A1(multiplier_0_n_12),.A2(multiplier_0_op2_reg[4]),.ZN(multiplier_0_n_26));
	NOR4_X1_LVT multiplier_0i_60_30 (.A1(multiplier_0_n_60_24),.A2(multiplier_0_n_60_25),.A3(multiplier_0_n_149),.A4(multiplier_0_n_26),.ZN(multiplier_0_n_60_26));
	AOI22_X1_LVT multiplier_0i_60_31 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[4]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[4]),.ZN(multiplier_0_n_60_27));
	OAI21_X1_LVT multiplier_0i_60_32 (.A(multiplier_0_n_60_26),.B1(multiplier_0_n_60_27),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[4]));
	AOI22_X1_LVT multiplier_0i_60_21 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_101),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_125),.ZN(multiplier_0_n_60_18));
	NOR2_X1_LVT multiplier_0i_60_22 (.A1(multiplier_0_n_60_18),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_19));
	AND2_X1_LVT multiplier_0i_60_23 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[3]),.ZN(multiplier_0_n_60_20));
	AND2_X1_LVT multiplier_0i_12_3 (.A1(multiplier_0_n_12),.A2(multiplier_0_op2_reg[3]),.ZN(multiplier_0_n_25));
	NOR4_X1_LVT multiplier_0i_60_24 (.A1(multiplier_0_n_60_19),.A2(multiplier_0_n_60_20),.A3(multiplier_0_n_149),.A4(multiplier_0_n_25),.ZN(multiplier_0_n_60_21));
	AOI22_X1_LVT multiplier_0i_60_25 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[3]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[3]),.ZN(multiplier_0_n_60_22));
	OAI21_X1_LVT multiplier_0i_60_26 (.A(multiplier_0_n_60_21),.B1(multiplier_0_n_60_22),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[3]));
	AOI22_X1_LVT multiplier_0i_60_15 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_102),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_124),.ZN(multiplier_0_n_60_13));
	NOR2_X1_LVT multiplier_0i_60_16 (.A1(multiplier_0_n_60_13),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_14));
	AND2_X1_LVT multiplier_0i_60_17 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[2]),.ZN(multiplier_0_n_60_15));
	AND2_X1_LVT multiplier_0i_12_2 (.A1(multiplier_0_n_12),.A2(multiplier_0_op2_reg[2]),.ZN(multiplier_0_n_24));
	NOR4_X1_LVT multiplier_0i_60_18 (.A1(multiplier_0_n_60_14),.A2(multiplier_0_n_60_15),.A3(multiplier_0_n_149),.A4(multiplier_0_n_24),.ZN(multiplier_0_n_60_16));
	AOI22_X1_LVT multiplier_0i_60_19 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[2]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[2]),.ZN(multiplier_0_n_60_17));
	OAI21_X1_LVT multiplier_0i_60_20 (.A(multiplier_0_n_60_16),.B1(multiplier_0_n_60_17),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[2]));
	AOI22_X1_LVT multiplier_0i_60_9 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_103),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_123),.ZN(multiplier_0_n_60_8));
	NOR2_X1_LVT multiplier_0i_60_10 (.A1(multiplier_0_n_60_8),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_9));
	AND2_X1_LVT multiplier_0i_60_11 (.A1(multiplier_0_n_150),.A2(multiplier_0_op1[1]),.ZN(multiplier_0_n_60_10));
	INV_X1_LVT multiplier_0i_55_0 (.A(multiplier_0_cycle[1]),.ZN(multiplier_0_n_55_0));
	AOI22_X1_LVT multiplier_0i_55_3 (.A1(multiplier_0_n_55_0),.A2(multiplier_0_sumext_s[1]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_sumext_s_nxt[1]),.ZN(multiplier_0_n_55_2));
	INV_X1_LVT multiplier_0i_55_4 (.A(multiplier_0_n_55_2),.ZN(multiplier_0_n_145));
	AND2_X1_LVT multiplier_0i_56_1 (.A1(multiplier_0_reg_rd15),.A2(multiplier_0_n_145),.ZN(multiplier_0_n_147));
	AND2_X1_LVT multiplier_0i_12_1 (.A1(multiplier_0_n_12),.A2(multiplier_0_op2_reg[1]),.ZN(multiplier_0_n_23));
	NOR4_X1_LVT multiplier_0i_60_12 (.A1(multiplier_0_n_60_9),.A2(multiplier_0_n_60_10),.A3(multiplier_0_n_147),.A4(multiplier_0_n_23),.ZN(multiplier_0_n_60_11));
	AOI22_X1_LVT multiplier_0i_60_13 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[1]),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_reshi_nxt[1]),.ZN(multiplier_0_n_60_12));
	OAI21_X1_LVT multiplier_0i_60_14 (.A(multiplier_0_n_60_11),.B1(multiplier_0_n_60_12),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[1]));
	AOI22_X1_LVT multiplier_0i_60_1 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_n_104),.B1(multiplier_0_cycle[1]),.B2(multiplier_0_n_122),.ZN(multiplier_0_n_60_1));
	NOR2_X1_LVT multiplier_0i_60_3 (.A1(multiplier_0_n_60_1),.A2(multiplier_0_n_60_2),.ZN(multiplier_0_n_60_3));
	AND2_X1_LVT multiplier_0i_60_4 (.A1(multiplier_0_op1[0]),.A2(multiplier_0_n_150),.ZN(multiplier_0_n_60_4));
	OR2_X1_LVT multiplier_0i_49_0 (.A1(multiplier_0_n_138),.A2(multiplier_0_sumext_s[0]),.ZN(multiplier_0_n_139));
	INV_X1_LVT multiplier_0i_50_1 (.A(multiplier_0_n_139),.ZN(multiplier_0_n_50_1));
	OAI21_X1_LVT multiplier_0i_50_2 (.A(multiplier_0_n_50_0),.B1(multiplier_0_n_50_1),.B2(multiplier_0_sign_sel),.ZN(multiplier_0_sumext_s_nxt[0]));
	AND2_X1_LVT multiplier_0i_52_1 (.A1(multiplier_0_n_52_0),.A2(multiplier_0_sumext_s_nxt[0]),.ZN(multiplier_0_n_141));
	DFFR_X1_LVT multiplier_0sumext_s_reg___05F05b0___05F05d (.D(multiplier_0_n_141),.RN(multiplier_0_n_38),.CK(multiplier_0_n_140),.Q(multiplier_0_sumext_s[0]),.QN());
	AOI22_X1_LVT multiplier_0i_55_1 (.A1(multiplier_0_n_55_0),.A2(multiplier_0_sumext_s[0]),.B1(multiplier_0_sumext_s_nxt[0]),.B2(multiplier_0_cycle[1]),.ZN(multiplier_0_n_55_1));
	INV_X1_LVT multiplier_0i_55_2 (.A(multiplier_0_n_55_1),.ZN(multiplier_0_n_144));
	AND2_X1_LVT multiplier_0i_56_0 (.A1(multiplier_0_n_144),.A2(multiplier_0_reg_rd15),.ZN(multiplier_0_n_146));
	AND2_X1_LVT multiplier_0i_12_0 (.A1(multiplier_0_op2_reg[0]),.A2(multiplier_0_n_12),.ZN(multiplier_0_n_22));
	NOR4_X1_LVT multiplier_0i_60_5 (.A1(multiplier_0_n_60_3),.A2(multiplier_0_n_60_4),.A3(multiplier_0_n_146),.A4(multiplier_0_n_22),.ZN(multiplier_0_n_60_5));
	AOI22_X1_LVT multiplier_0i_60_6 (.A1(multiplier_0_n_60_0),.A2(multiplier_0_reshi[0]),.B1(multiplier_0_reshi_nxt[0]),.B2(multiplier_0_cycle[1]),.ZN(multiplier_0_n_60_6));
	OAI21_X1_LVT multiplier_0i_60_8 (.A(multiplier_0_n_60_5),.B1(multiplier_0_n_60_6),.B2(multiplier_0_n_60_7),.ZN(per_dout_mpy[0]));
	OR4_X1_LVT i_0_0_30 (.A1(per_dout_mpy[15]),.A2(per_dout_wdog[15]),.A3(per_dout_sfr[15]),.A4(per_dout_clk[15]),.ZN(n_0_0_15));
	OR2_X1_LVT i_0_0_31 (.A1(n_0_0_15),.A2(per_dout[15]),.ZN(per_dout_or[15]));
	OR4_X1_LVT i_0_0_28 (.A1(per_dout_mpy[14]),.A2(per_dout_wdog[14]),.A3(per_dout_sfr[14]),.A4(per_dout_clk[14]),.ZN(n_0_0_14));
	OR2_X1_LVT i_0_0_29 (.A1(n_0_0_14),.A2(per_dout[14]),.ZN(per_dout_or[14]));
	OR4_X1_LVT i_0_0_26 (.A1(per_dout_mpy[13]),.A2(per_dout_wdog[13]),.A3(per_dout_sfr[13]),.A4(per_dout_clk[13]),.ZN(n_0_0_13));
	OR2_X1_LVT i_0_0_27 (.A1(n_0_0_13),.A2(per_dout[13]),.ZN(per_dout_or[13]));
	OR4_X1_LVT i_0_0_24 (.A1(per_dout_mpy[12]),.A2(per_dout_wdog[12]),.A3(per_dout_sfr[12]),.A4(per_dout_clk[12]),.ZN(n_0_0_12));
	OR2_X1_LVT i_0_0_25 (.A1(n_0_0_12),.A2(per_dout[12]),.ZN(per_dout_or[12]));
	OR4_X1_LVT i_0_0_22 (.A1(per_dout_mpy[11]),.A2(per_dout_wdog[11]),.A3(per_dout_sfr[11]),.A4(per_dout_clk[11]),.ZN(n_0_0_11));
	OR2_X1_LVT i_0_0_23 (.A1(n_0_0_11),.A2(per_dout[11]),.ZN(per_dout_or[11]));
	OR4_X1_LVT i_0_0_20 (.A1(per_dout_mpy[10]),.A2(per_dout_wdog[10]),.A3(per_dout_sfr[10]),.A4(per_dout_clk[10]),.ZN(n_0_0_10));
	OR2_X1_LVT i_0_0_21 (.A1(n_0_0_10),.A2(per_dout[10]),.ZN(per_dout_or[10]));
	OR4_X1_LVT i_0_0_18 (.A1(per_dout_mpy[9]),.A2(per_dout_wdog[9]),.A3(per_dout_sfr[9]),.A4(per_dout_clk[9]),.ZN(n_0_0_9));
	OR2_X1_LVT i_0_0_19 (.A1(n_0_0_9),.A2(per_dout[9]),.ZN(per_dout_or[9]));
	OR4_X1_LVT i_0_0_16 (.A1(per_dout_mpy[8]),.A2(per_dout_wdog[8]),.A3(per_dout_sfr[8]),.A4(per_dout_clk[8]),.ZN(n_0_0_8));
	OR2_X1_LVT i_0_0_17 (.A1(n_0_0_8),.A2(per_dout[8]),.ZN(per_dout_or[8]));
	OR4_X1_LVT i_0_0_14 (.A1(per_dout_mpy[7]),.A2(per_dout_wdog[7]),.A3(per_dout_sfr[7]),.A4(per_dout_clk[7]),.ZN(n_0_0_7));
	OR2_X1_LVT i_0_0_15 (.A1(n_0_0_7),.A2(per_dout[7]),.ZN(per_dout_or[7]));
	OR4_X1_LVT i_0_0_12 (.A1(per_dout_mpy[6]),.A2(per_dout_wdog[6]),.A3(per_dout_sfr[6]),.A4(per_dout_clk[6]),.ZN(n_0_0_6));
	OR2_X1_LVT i_0_0_13 (.A1(n_0_0_6),.A2(per_dout[6]),.ZN(per_dout_or[6]));
	OR4_X1_LVT i_0_0_10 (.A1(per_dout_mpy[5]),.A2(per_dout_wdog[5]),.A3(per_dout_sfr[5]),.A4(per_dout_clk[5]),.ZN(n_0_0_5));
	OR2_X1_LVT i_0_0_11 (.A1(n_0_0_5),.A2(per_dout[5]),.ZN(per_dout_or[5]));
	OR4_X1_LVT i_0_0_8 (.A1(per_dout_mpy[4]),.A2(per_dout_wdog[4]),.A3(per_dout_sfr[4]),.A4(per_dout_clk[4]),.ZN(n_0_0_4));
	OR2_X1_LVT i_0_0_9 (.A1(n_0_0_4),.A2(per_dout[4]),.ZN(per_dout_or[4]));
	OR4_X1_LVT i_0_0_6 (.A1(per_dout_mpy[3]),.A2(per_dout_wdog[3]),.A3(per_dout_sfr[3]),.A4(per_dout_clk[3]),.ZN(n_0_0_3));
	OR2_X1_LVT i_0_0_7 (.A1(n_0_0_3),.A2(per_dout[3]),.ZN(per_dout_or[3]));
	OR4_X1_LVT i_0_0_4 (.A1(per_dout_mpy[2]),.A2(per_dout_wdog[2]),.A3(per_dout_sfr[2]),.A4(per_dout_clk[2]),.ZN(n_0_0_2));
	OR2_X1_LVT i_0_0_5 (.A1(n_0_0_2),.A2(per_dout[2]),.ZN(per_dout_or[2]));
	OR4_X1_LVT i_0_0_2 (.A1(per_dout_mpy[1]),.A2(per_dout_wdog[1]),.A3(per_dout_sfr[1]),.A4(per_dout_clk[1]),.ZN(n_0_0_1));
	OR2_X1_LVT i_0_0_3 (.A1(n_0_0_1),.A2(per_dout[1]),.ZN(per_dout_or[1]));
	OR4_X1_LVT i_0_0_0 (.A1(per_dout_mpy[0]),.A2(per_dout_wdog[0]),.A3(per_dout_sfr[0]),.A4(per_dout_clk[0]),.ZN(n_0_0_0));
	OR2_X1_LVT i_0_0_1 (.A1(n_0_0_0),.A2(per_dout[0]),.ZN(per_dout_or[0]));
	AOI21_X1_LVT mem_backbone_0i_0_0 (.A(dbg_halt_cmd),.B1(dma_en),.B2(dma_priority),.ZN(mem_backbone_0_n_0_0));
	INV_X1_LVT mem_backbone_0i_0_1 (.A(mem_backbone_0_n_0_0),.ZN(cpu_halt_cmd));
	OR2_X1_LVT mem_backbone_0i_4_0 (.A1(dbg_mem_en),.A2(dma_en),.ZN(mem_backbone_0_ext_mem_en));
	AND4_X1_LVT mem_backbone_0i_8_0 (.A1(n_2),.A2(n_1),.A3(n_0),.A4(fe_mb_en),.ZN(mem_backbone_0_n_8_0));
	AND2_X1_LVT mem_backbone_0i_8_1 (.A1(mem_backbone_0_n_8_0),.A2(n_3),.ZN(mem_backbone_0_fe_pmem_en));
	INV_X1_LVT mem_backbone_0i_9_0 (.A(mem_backbone_0_fe_pmem_en),.ZN(mem_backbone_0_n_0));
	INV_X1_LVT mem_backbone_0i_2_0 (.A(dbg_mem_en),.ZN(mem_backbone_0_n_2_0));
	AOI22_X1_LVT mem_backbone_0i_2_23 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[11]),.B1(dbg_mem_en),.B2(dbg_mem_addr[12]),.ZN(mem_backbone_0_n_2_12));
	INV_X1_LVT mem_backbone_0i_2_24 (.A(mem_backbone_0_n_2_12),.ZN(mem_backbone_0_ext_mem_addr[11]));
	AOI22_X1_LVT mem_backbone_0i_2_25 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[12]),.B1(dbg_mem_en),.B2(dbg_mem_addr[13]),.ZN(mem_backbone_0_n_2_13));
	INV_X1_LVT mem_backbone_0i_2_26 (.A(mem_backbone_0_n_2_13),.ZN(mem_backbone_0_ext_mem_addr[12]));
	AOI22_X1_LVT mem_backbone_0i_2_27 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[13]),.B1(dbg_mem_en),.B2(dbg_mem_addr[14]),.ZN(mem_backbone_0_n_2_14));
	INV_X1_LVT mem_backbone_0i_2_28 (.A(mem_backbone_0_n_2_14),.ZN(mem_backbone_0_ext_mem_addr[13]));
	AOI22_X1_LVT mem_backbone_0i_2_29 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[14]),.B1(dbg_mem_en),.B2(dbg_mem_addr[15]),.ZN(mem_backbone_0_n_2_15));
	INV_X1_LVT mem_backbone_0i_2_30 (.A(mem_backbone_0_n_2_15),.ZN(mem_backbone_0_ext_mem_addr[14]));
	AND4_X1_LVT mem_backbone_0i_7_0 (.A1(mem_backbone_0_ext_mem_addr[11]),.A2(mem_backbone_0_ext_mem_addr[12]),.A3(mem_backbone_0_ext_mem_addr[13]),.A4(mem_backbone_0_ext_mem_addr[14]),.ZN(mem_backbone_0_ext_pmem_sel));
	NAND3_X1_LVT mem_backbone_0i_12_0 (.A1(mem_backbone_0_ext_mem_en),.A2(mem_backbone_0_n_0),.A3(mem_backbone_0_ext_pmem_sel),.ZN(mem_backbone_0_n_12_0));
	NOR2_X1_LVT mem_backbone_0i_10_0 (.A1(eu_mb_wr[0]),.A2(eu_mb_wr[1]),.ZN(mem_backbone_0_n_1));
	NAND4_X1_LVT mem_backbone_0i_11_0 (.A1(eu_mab[14]),.A2(eu_mab[15]),.A3(eu_mb_en),.A4(mem_backbone_0_n_1),.ZN(mem_backbone_0_n_11_0));
	NAND2_X1_LVT mem_backbone_0i_11_1 (.A1(eu_mab[12]),.A2(eu_mab[13]),.ZN(mem_backbone_0_n_11_1));
	NOR2_X1_LVT mem_backbone_0i_11_2 (.A1(mem_backbone_0_n_11_0),.A2(mem_backbone_0_n_11_1),.ZN(mem_backbone_0_eu_pmem_en));
	NOR2_X1_LVT mem_backbone_0i_12_1 (.A1(mem_backbone_0_n_12_0),.A2(mem_backbone_0_eu_pmem_en),.ZN(mem_backbone_0_ext_pmem_en));
	INV_X1_LVT mem_backbone_0i_13_0 (.A(puc_rst),.ZN(mem_backbone_0_n_2));
	DFFR_X1_LVT mem_backbone_0ext_mem_din_sel_reg___05F05b1___05F05d (.D(mem_backbone_0_ext_pmem_en),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_ext_mem_din_sel[1]),.QN());
	OR4_X1_LVT mem_backbone_0i_3_0 (.A1(mem_backbone_0_ext_mem_addr[11]),.A2(mem_backbone_0_ext_mem_addr[12]),.A3(mem_backbone_0_ext_mem_addr[13]),.A4(mem_backbone_0_ext_mem_addr[14]),.ZN(mem_backbone_0_n_3_0));
	AOI22_X1_LVT mem_backbone_0i_2_17 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[8]),.B1(dbg_mem_en),.B2(dbg_mem_addr[9]),.ZN(mem_backbone_0_n_2_9));
	INV_X1_LVT mem_backbone_0i_2_18 (.A(mem_backbone_0_n_2_9),.ZN(mem_backbone_0_ext_mem_addr[8]));
	AOI22_X1_LVT mem_backbone_0i_2_19 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[9]),.B1(dbg_mem_en),.B2(dbg_mem_addr[10]),.ZN(mem_backbone_0_n_2_10));
	INV_X1_LVT mem_backbone_0i_2_20 (.A(mem_backbone_0_n_2_10),.ZN(mem_backbone_0_ext_mem_addr[9]));
	AOI22_X1_LVT mem_backbone_0i_2_21 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[10]),.B1(dbg_mem_en),.B2(dbg_mem_addr[11]),.ZN(mem_backbone_0_n_2_11));
	INV_X1_LVT mem_backbone_0i_2_22 (.A(mem_backbone_0_n_2_11),.ZN(mem_backbone_0_ext_mem_addr[10]));
	NOR4_X1_LVT mem_backbone_0i_3_1 (.A1(mem_backbone_0_n_3_0),.A2(mem_backbone_0_ext_mem_addr[8]),.A3(mem_backbone_0_ext_mem_addr[9]),.A4(mem_backbone_0_ext_mem_addr[10]),.ZN(mem_backbone_0_ext_per_sel));
	NAND2_X1_LVT mem_backbone_0i_6_0 (.A1(mem_backbone_0_ext_mem_en),.A2(mem_backbone_0_ext_per_sel),.ZN(mem_backbone_0_n_6_0));
	INV_X1_LVT mem_backbone_0i_5_0 (.A(eu_mb_en),.ZN(mem_backbone_0_n_5_0));
	NOR4_X1_LVT mem_backbone_0i_5_1 (.A1(mem_backbone_0_n_5_0),.A2(eu_mab[13]),.A3(eu_mab[14]),.A4(eu_mab[15]),.ZN(mem_backbone_0_n_5_1));
	NOR4_X1_LVT mem_backbone_0i_5_2 (.A1(eu_mab[9]),.A2(eu_mab[10]),.A3(eu_mab[11]),.A4(eu_mab[12]),.ZN(mem_backbone_0_n_5_2));
	AND2_X1_LVT mem_backbone_0i_5_3 (.A1(mem_backbone_0_n_5_1),.A2(mem_backbone_0_n_5_2),.ZN(mem_backbone_0_eu_per_en));
	NOR2_X1_LVT mem_backbone_0i_6_1 (.A1(mem_backbone_0_n_6_0),.A2(mem_backbone_0_eu_per_en),.ZN(mem_backbone_0_ext_per_en));
	DFFR_X1_LVT mem_backbone_0ext_mem_din_sel_reg___05F05b0___05F05d (.D(mem_backbone_0_ext_per_en),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_ext_mem_din_sel[0]),.QN());
	INV_X1_LVT mem_backbone_0i_15_1 (.A(mem_backbone_0_ext_mem_din_sel[0]),.ZN(mem_backbone_0_n_15_0));
	NOR2_X1_LVT mem_backbone_0i_15_2 (.A1(mem_backbone_0_n_15_0),.A2(mem_backbone_0_ext_mem_din_sel[1]),.ZN(mem_backbone_0_n_4));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b15___05F05d (.D(per_dout_or[15]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[15]),.QN());
	NOR2_X1_LVT mem_backbone_0i_15_0 (.A1(mem_backbone_0_ext_mem_din_sel[0]),.A2(mem_backbone_0_ext_mem_din_sel[1]),.ZN(mem_backbone_0_n_3));
	AOI222_X1_LVT mem_backbone_0i_16_30 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[15]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[15]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[15]),.ZN(mem_backbone_0_n_16_15));
	INV_X1_LVT mem_backbone_0i_16_31 (.A(mem_backbone_0_n_16_15),.ZN(dbg_mem_din[15]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b14___05F05d (.D(per_dout_or[14]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[14]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_28 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[14]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[14]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[14]),.ZN(mem_backbone_0_n_16_14));
	INV_X1_LVT mem_backbone_0i_16_29 (.A(mem_backbone_0_n_16_14),.ZN(dbg_mem_din[14]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b13___05F05d (.D(per_dout_or[13]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[13]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_26 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[13]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[13]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[13]),.ZN(mem_backbone_0_n_16_13));
	INV_X1_LVT mem_backbone_0i_16_27 (.A(mem_backbone_0_n_16_13),.ZN(dbg_mem_din[13]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b12___05F05d (.D(per_dout_or[12]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[12]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_24 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[12]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[12]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[12]),.ZN(mem_backbone_0_n_16_12));
	INV_X1_LVT mem_backbone_0i_16_25 (.A(mem_backbone_0_n_16_12),.ZN(dbg_mem_din[12]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b11___05F05d (.D(per_dout_or[11]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[11]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_22 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[11]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[11]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[11]),.ZN(mem_backbone_0_n_16_11));
	INV_X1_LVT mem_backbone_0i_16_23 (.A(mem_backbone_0_n_16_11),.ZN(dbg_mem_din[11]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b10___05F05d (.D(per_dout_or[10]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[10]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_20 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[10]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[10]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[10]),.ZN(mem_backbone_0_n_16_10));
	INV_X1_LVT mem_backbone_0i_16_21 (.A(mem_backbone_0_n_16_10),.ZN(dbg_mem_din[10]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b9___05F05d (.D(per_dout_or[9]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[9]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_18 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[9]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[9]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[9]),.ZN(mem_backbone_0_n_16_9));
	INV_X1_LVT mem_backbone_0i_16_19 (.A(mem_backbone_0_n_16_9),.ZN(dbg_mem_din[9]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b8___05F05d (.D(per_dout_or[8]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[8]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_16 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[8]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[8]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[8]),.ZN(mem_backbone_0_n_16_8));
	INV_X1_LVT mem_backbone_0i_16_17 (.A(mem_backbone_0_n_16_8),.ZN(dbg_mem_din[8]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b7___05F05d (.D(per_dout_or[7]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[7]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_14 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[7]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[7]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[7]),.ZN(mem_backbone_0_n_16_7));
	INV_X1_LVT mem_backbone_0i_16_15 (.A(mem_backbone_0_n_16_7),.ZN(dbg_mem_din[7]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b6___05F05d (.D(per_dout_or[6]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[6]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_12 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[6]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[6]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[6]),.ZN(mem_backbone_0_n_16_6));
	INV_X1_LVT mem_backbone_0i_16_13 (.A(mem_backbone_0_n_16_6),.ZN(dbg_mem_din[6]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b5___05F05d (.D(per_dout_or[5]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[5]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_10 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[5]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[5]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[5]),.ZN(mem_backbone_0_n_16_5));
	INV_X1_LVT mem_backbone_0i_16_11 (.A(mem_backbone_0_n_16_5),.ZN(dbg_mem_din[5]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b4___05F05d (.D(per_dout_or[4]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[4]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_8 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[4]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[4]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[4]),.ZN(mem_backbone_0_n_16_4));
	INV_X1_LVT mem_backbone_0i_16_9 (.A(mem_backbone_0_n_16_4),.ZN(dbg_mem_din[4]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b3___05F05d (.D(per_dout_or[3]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[3]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_6 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[3]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[3]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[3]),.ZN(mem_backbone_0_n_16_3));
	INV_X1_LVT mem_backbone_0i_16_7 (.A(mem_backbone_0_n_16_3),.ZN(dbg_mem_din[3]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b2___05F05d (.D(per_dout_or[2]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[2]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_4 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[2]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[2]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[2]),.ZN(mem_backbone_0_n_16_2));
	INV_X1_LVT mem_backbone_0i_16_5 (.A(mem_backbone_0_n_16_2),.ZN(dbg_mem_din[2]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b1___05F05d (.D(per_dout_or[1]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[1]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_2 (.A1(mem_backbone_0_ext_mem_din_sel[1]),.A2(pmem_dout[1]),.B1(mem_backbone_0_n_4),.B2(mem_backbone_0_per_dout_val[1]),.C1(mem_backbone_0_n_3),.C2(dmem_dout[1]),.ZN(mem_backbone_0_n_16_1));
	INV_X1_LVT mem_backbone_0i_16_3 (.A(mem_backbone_0_n_16_1),.ZN(dbg_mem_din[1]));
	DFFR_X1_LVT mem_backbone_0per_dout_val_reg___05F05b0___05F05d (.D(per_dout_or[0]),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_per_dout_val[0]),.QN());
	AOI222_X1_LVT mem_backbone_0i_16_0 (.A1(pmem_dout[0]),.A2(mem_backbone_0_ext_mem_din_sel[1]),.B1(mem_backbone_0_per_dout_val[0]),.B2(mem_backbone_0_n_4),.C1(dmem_dout[0]),.C2(mem_backbone_0_n_3),.ZN(mem_backbone_0_n_16_0));
	INV_X1_LVT mem_backbone_0i_16_1 (.A(mem_backbone_0_n_16_0),.ZN(dbg_mem_din[0]));
	INV_X1_LVT mem_backbone_0i_19_0 (.A(mem_backbone_0_ext_mem_addr[11]),.ZN(mem_backbone_0_n_19_0));
	INV_X1_LVT mem_backbone_0i_19_1 (.A(mem_backbone_0_ext_mem_addr[12]),.ZN(mem_backbone_0_n_19_1));
	INV_X1_LVT mem_backbone_0i_19_2 (.A(mem_backbone_0_ext_mem_addr[13]),.ZN(mem_backbone_0_n_19_2));
	INV_X1_LVT mem_backbone_0i_19_3 (.A(mem_backbone_0_ext_mem_addr[14]),.ZN(mem_backbone_0_n_19_3));
	NAND4_X1_LVT mem_backbone_0i_19_4 (.A1(mem_backbone_0_n_19_0),.A2(mem_backbone_0_n_19_1),.A3(mem_backbone_0_n_19_2),.A4(mem_backbone_0_n_19_3),.ZN(mem_backbone_0_n_19_4));
	NOR4_X1_LVT mem_backbone_0i_19_5 (.A1(mem_backbone_0_n_19_4),.A2(mem_backbone_0_ext_mem_addr[8]),.A3(mem_backbone_0_ext_mem_addr[9]),.A4(mem_backbone_0_ext_mem_addr[10]),.ZN(mem_backbone_0_n_19_5));
	AND2_X1_LVT mem_backbone_0i_19_6 (.A1(mem_backbone_0_ext_mem_addr[8]),.A2(mem_backbone_0_ext_mem_addr[9]),.ZN(mem_backbone_0_n_19_6));
	NOR4_X1_LVT mem_backbone_0i_19_7 (.A1(mem_backbone_0_n_19_4),.A2(mem_backbone_0_n_19_5),.A3(mem_backbone_0_n_19_6),.A4(mem_backbone_0_ext_mem_addr[10]),.ZN(mem_backbone_0_ext_dmem_sel));
	NAND2_X1_LVT mem_backbone_0i_21_0 (.A1(mem_backbone_0_ext_mem_en),.A2(mem_backbone_0_ext_dmem_sel),.ZN(mem_backbone_0_n_21_0));
	OR4_X1_LVT mem_backbone_0i_20_0 (.A1(eu_mab[12]),.A2(eu_mab[13]),.A3(eu_mab[14]),.A4(eu_mab[15]),.ZN(mem_backbone_0_n_20_0));
	NOR4_X1_LVT mem_backbone_0i_20_1 (.A1(mem_backbone_0_n_20_0),.A2(eu_mab[9]),.A3(eu_mab[10]),.A4(eu_mab[11]),.ZN(mem_backbone_0_n_20_1));
	AND2_X1_LVT mem_backbone_0i_20_2 (.A1(eu_mab[9]),.A2(eu_mab[10]),.ZN(mem_backbone_0_n_20_2));
	NOR4_X1_LVT mem_backbone_0i_20_3 (.A1(mem_backbone_0_n_20_1),.A2(mem_backbone_0_n_20_2),.A3(eu_mab[11]),.A4(eu_mab[12]),.ZN(mem_backbone_0_n_20_3));
	INV_X1_LVT mem_backbone_0i_20_4 (.A(eu_mb_en),.ZN(mem_backbone_0_n_20_4));
	NOR4_X1_LVT mem_backbone_0i_20_5 (.A1(mem_backbone_0_n_20_4),.A2(eu_mab[13]),.A3(eu_mab[14]),.A4(eu_mab[15]),.ZN(mem_backbone_0_n_20_5));
	AND2_X1_LVT mem_backbone_0i_20_6 (.A1(mem_backbone_0_n_20_3),.A2(mem_backbone_0_n_20_5),.ZN(mem_backbone_0_eu_dmem_en));
	NOR2_X1_LVT mem_backbone_0i_21_1 (.A1(mem_backbone_0_n_21_0),.A2(mem_backbone_0_eu_dmem_en),.ZN(mem_backbone_0_ext_dmem_en));
	INV_X1_LVT mem_backbone_0i_22_0 (.A(mem_backbone_0_ext_dmem_en),.ZN(mem_backbone_0_n_22_0));
	INV_X1_LVT mem_backbone_0i_17_0 (.A(eu_mab[9]),.ZN(mem_backbone_0_n_5));
	INV_X1_LVT mem_backbone_0i_18_0 (.A(mem_backbone_0_ext_mem_addr[8]),.ZN(mem_backbone_0_n_6));
	AOI22_X1_LVT mem_backbone_0i_22_17 (.A1(mem_backbone_0_n_22_0),.A2(mem_backbone_0_n_5),.B1(mem_backbone_0_ext_dmem_en),.B2(mem_backbone_0_n_6),.ZN(mem_backbone_0_n_22_9));
	INV_X1_LVT mem_backbone_0i_22_18 (.A(mem_backbone_0_n_22_9),.ZN(dmem_addr[8]));
	AOI22_X1_LVT mem_backbone_0i_2_15 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[7]),.B1(dbg_mem_en),.B2(dbg_mem_addr[8]),.ZN(mem_backbone_0_n_2_8));
	INV_X1_LVT mem_backbone_0i_2_16 (.A(mem_backbone_0_n_2_8),.ZN(mem_backbone_0_ext_mem_addr[7]));
	AOI22_X1_LVT mem_backbone_0i_22_15 (.A1(mem_backbone_0_n_22_0),.A2(eu_mab[8]),.B1(mem_backbone_0_ext_dmem_en),.B2(mem_backbone_0_ext_mem_addr[7]),.ZN(mem_backbone_0_n_22_8));
	INV_X1_LVT mem_backbone_0i_22_16 (.A(mem_backbone_0_n_22_8),.ZN(dmem_addr[7]));
	AOI22_X1_LVT mem_backbone_0i_2_13 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[6]),.B1(dbg_mem_en),.B2(dbg_mem_addr[7]),.ZN(mem_backbone_0_n_2_7));
	INV_X1_LVT mem_backbone_0i_2_14 (.A(mem_backbone_0_n_2_7),.ZN(mem_backbone_0_ext_mem_addr[6]));
	AOI22_X1_LVT mem_backbone_0i_22_13 (.A1(mem_backbone_0_n_22_0),.A2(eu_mab[7]),.B1(mem_backbone_0_ext_dmem_en),.B2(mem_backbone_0_ext_mem_addr[6]),.ZN(mem_backbone_0_n_22_7));
	INV_X1_LVT mem_backbone_0i_22_14 (.A(mem_backbone_0_n_22_7),.ZN(dmem_addr[6]));
	AOI22_X1_LVT mem_backbone_0i_2_11 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[5]),.B1(dbg_mem_en),.B2(dbg_mem_addr[6]),.ZN(mem_backbone_0_n_2_6));
	INV_X1_LVT mem_backbone_0i_2_12 (.A(mem_backbone_0_n_2_6),.ZN(mem_backbone_0_ext_mem_addr[5]));
	AOI22_X1_LVT mem_backbone_0i_22_11 (.A1(mem_backbone_0_n_22_0),.A2(eu_mab[6]),.B1(mem_backbone_0_ext_dmem_en),.B2(mem_backbone_0_ext_mem_addr[5]),.ZN(mem_backbone_0_n_22_6));
	INV_X1_LVT mem_backbone_0i_22_12 (.A(mem_backbone_0_n_22_6),.ZN(dmem_addr[5]));
	AOI22_X1_LVT mem_backbone_0i_2_9 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[4]),.B1(dbg_mem_en),.B2(dbg_mem_addr[5]),.ZN(mem_backbone_0_n_2_5));
	INV_X1_LVT mem_backbone_0i_2_10 (.A(mem_backbone_0_n_2_5),.ZN(mem_backbone_0_ext_mem_addr[4]));
	AOI22_X1_LVT mem_backbone_0i_22_9 (.A1(mem_backbone_0_n_22_0),.A2(eu_mab[5]),.B1(mem_backbone_0_ext_dmem_en),.B2(mem_backbone_0_ext_mem_addr[4]),.ZN(mem_backbone_0_n_22_5));
	INV_X1_LVT mem_backbone_0i_22_10 (.A(mem_backbone_0_n_22_5),.ZN(dmem_addr[4]));
	AOI22_X1_LVT mem_backbone_0i_2_7 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[3]),.B1(dbg_mem_en),.B2(dbg_mem_addr[4]),.ZN(mem_backbone_0_n_2_4));
	INV_X1_LVT mem_backbone_0i_2_8 (.A(mem_backbone_0_n_2_4),.ZN(mem_backbone_0_ext_mem_addr[3]));
	AOI22_X1_LVT mem_backbone_0i_22_7 (.A1(mem_backbone_0_n_22_0),.A2(eu_mab[4]),.B1(mem_backbone_0_ext_dmem_en),.B2(mem_backbone_0_ext_mem_addr[3]),.ZN(mem_backbone_0_n_22_4));
	INV_X1_LVT mem_backbone_0i_22_8 (.A(mem_backbone_0_n_22_4),.ZN(dmem_addr[3]));
	AOI22_X1_LVT mem_backbone_0i_2_5 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[2]),.B1(dbg_mem_en),.B2(dbg_mem_addr[3]),.ZN(mem_backbone_0_n_2_3));
	INV_X1_LVT mem_backbone_0i_2_6 (.A(mem_backbone_0_n_2_3),.ZN(mem_backbone_0_ext_mem_addr[2]));
	AOI22_X1_LVT mem_backbone_0i_22_5 (.A1(mem_backbone_0_n_22_0),.A2(eu_mab[3]),.B1(mem_backbone_0_ext_dmem_en),.B2(mem_backbone_0_ext_mem_addr[2]),.ZN(mem_backbone_0_n_22_3));
	INV_X1_LVT mem_backbone_0i_22_6 (.A(mem_backbone_0_n_22_3),.ZN(dmem_addr[2]));
	AOI22_X1_LVT mem_backbone_0i_2_3 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[1]),.B1(dbg_mem_en),.B2(dbg_mem_addr[2]),.ZN(mem_backbone_0_n_2_2));
	INV_X1_LVT mem_backbone_0i_2_4 (.A(mem_backbone_0_n_2_2),.ZN(mem_backbone_0_ext_mem_addr[1]));
	AOI22_X1_LVT mem_backbone_0i_22_3 (.A1(mem_backbone_0_n_22_0),.A2(eu_mab[2]),.B1(mem_backbone_0_ext_dmem_en),.B2(mem_backbone_0_ext_mem_addr[1]),.ZN(mem_backbone_0_n_22_2));
	INV_X1_LVT mem_backbone_0i_22_4 (.A(mem_backbone_0_n_22_2),.ZN(dmem_addr[1]));
	AOI22_X1_LVT mem_backbone_0i_2_1 (.A1(mem_backbone_0_n_2_0),.A2(dma_addr[0]),.B1(dbg_mem_addr[1]),.B2(dbg_mem_en),.ZN(mem_backbone_0_n_2_1));
	INV_X1_LVT mem_backbone_0i_2_2 (.A(mem_backbone_0_n_2_1),.ZN(mem_backbone_0_ext_mem_addr[0]));
	AOI22_X1_LVT mem_backbone_0i_22_1 (.A1(mem_backbone_0_n_22_0),.A2(eu_mab[1]),.B1(mem_backbone_0_ext_mem_addr[0]),.B2(mem_backbone_0_ext_dmem_en),.ZN(mem_backbone_0_n_22_1));
	INV_X1_LVT mem_backbone_0i_22_2 (.A(mem_backbone_0_n_22_1),.ZN(dmem_addr[0]));
	NOR2_X1_LVT mem_backbone_0i_23_0 (.A1(mem_backbone_0_ext_dmem_en),.A2(mem_backbone_0_eu_dmem_en),.ZN(dmem_cen));
	INV_X1_LVT mem_backbone_0i_25_0 (.A(mem_backbone_0_ext_dmem_en),.ZN(mem_backbone_0_n_25_0));
	INV_X1_LVT mem_backbone_0i_24_0 (.A(dbg_mem_en),.ZN(mem_backbone_0_n_24_0));
	AOI22_X1_LVT mem_backbone_0i_24_31 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[15]),.B1(dbg_mem_en),.B2(dbg_mem_dout[15]),.ZN(mem_backbone_0_n_24_16));
	INV_X1_LVT mem_backbone_0i_24_32 (.A(mem_backbone_0_n_24_16),.ZN(pmem_din[15]));
	AOI22_X1_LVT mem_backbone_0i_25_31 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[15]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[15]),.ZN(mem_backbone_0_n_25_16));
	INV_X1_LVT mem_backbone_0i_25_32 (.A(mem_backbone_0_n_25_16),.ZN(dmem_din[15]));
	AOI22_X1_LVT mem_backbone_0i_24_29 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[14]),.B1(dbg_mem_en),.B2(dbg_mem_dout[14]),.ZN(mem_backbone_0_n_24_15));
	INV_X1_LVT mem_backbone_0i_24_30 (.A(mem_backbone_0_n_24_15),.ZN(pmem_din[14]));
	AOI22_X1_LVT mem_backbone_0i_25_29 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[14]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[14]),.ZN(mem_backbone_0_n_25_15));
	INV_X1_LVT mem_backbone_0i_25_30 (.A(mem_backbone_0_n_25_15),.ZN(dmem_din[14]));
	AOI22_X1_LVT mem_backbone_0i_24_27 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[13]),.B1(dbg_mem_en),.B2(dbg_mem_dout[13]),.ZN(mem_backbone_0_n_24_14));
	INV_X1_LVT mem_backbone_0i_24_28 (.A(mem_backbone_0_n_24_14),.ZN(pmem_din[13]));
	AOI22_X1_LVT mem_backbone_0i_25_27 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[13]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[13]),.ZN(mem_backbone_0_n_25_14));
	INV_X1_LVT mem_backbone_0i_25_28 (.A(mem_backbone_0_n_25_14),.ZN(dmem_din[13]));
	AOI22_X1_LVT mem_backbone_0i_24_25 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[12]),.B1(dbg_mem_en),.B2(dbg_mem_dout[12]),.ZN(mem_backbone_0_n_24_13));
	INV_X1_LVT mem_backbone_0i_24_26 (.A(mem_backbone_0_n_24_13),.ZN(pmem_din[12]));
	AOI22_X1_LVT mem_backbone_0i_25_25 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[12]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[12]),.ZN(mem_backbone_0_n_25_13));
	INV_X1_LVT mem_backbone_0i_25_26 (.A(mem_backbone_0_n_25_13),.ZN(dmem_din[12]));
	AOI22_X1_LVT mem_backbone_0i_24_23 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[11]),.B1(dbg_mem_en),.B2(dbg_mem_dout[11]),.ZN(mem_backbone_0_n_24_12));
	INV_X1_LVT mem_backbone_0i_24_24 (.A(mem_backbone_0_n_24_12),.ZN(pmem_din[11]));
	AOI22_X1_LVT mem_backbone_0i_25_23 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[11]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[11]),.ZN(mem_backbone_0_n_25_12));
	INV_X1_LVT mem_backbone_0i_25_24 (.A(mem_backbone_0_n_25_12),.ZN(dmem_din[11]));
	AOI22_X1_LVT mem_backbone_0i_24_21 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[10]),.B1(dbg_mem_en),.B2(dbg_mem_dout[10]),.ZN(mem_backbone_0_n_24_11));
	INV_X1_LVT mem_backbone_0i_24_22 (.A(mem_backbone_0_n_24_11),.ZN(pmem_din[10]));
	AOI22_X1_LVT mem_backbone_0i_25_21 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[10]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[10]),.ZN(mem_backbone_0_n_25_11));
	INV_X1_LVT mem_backbone_0i_25_22 (.A(mem_backbone_0_n_25_11),.ZN(dmem_din[10]));
	AOI22_X1_LVT mem_backbone_0i_24_19 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[9]),.B1(dbg_mem_en),.B2(dbg_mem_dout[9]),.ZN(mem_backbone_0_n_24_10));
	INV_X1_LVT mem_backbone_0i_24_20 (.A(mem_backbone_0_n_24_10),.ZN(pmem_din[9]));
	AOI22_X1_LVT mem_backbone_0i_25_19 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[9]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[9]),.ZN(mem_backbone_0_n_25_10));
	INV_X1_LVT mem_backbone_0i_25_20 (.A(mem_backbone_0_n_25_10),.ZN(dmem_din[9]));
	AOI22_X1_LVT mem_backbone_0i_24_17 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[8]),.B1(dbg_mem_en),.B2(dbg_mem_dout[8]),.ZN(mem_backbone_0_n_24_9));
	INV_X1_LVT mem_backbone_0i_24_18 (.A(mem_backbone_0_n_24_9),.ZN(pmem_din[8]));
	AOI22_X1_LVT mem_backbone_0i_25_17 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[8]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[8]),.ZN(mem_backbone_0_n_25_9));
	INV_X1_LVT mem_backbone_0i_25_18 (.A(mem_backbone_0_n_25_9),.ZN(dmem_din[8]));
	AOI22_X1_LVT mem_backbone_0i_24_15 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[7]),.B1(dbg_mem_en),.B2(dbg_mem_dout[7]),.ZN(mem_backbone_0_n_24_8));
	INV_X1_LVT mem_backbone_0i_24_16 (.A(mem_backbone_0_n_24_8),.ZN(pmem_din[7]));
	AOI22_X1_LVT mem_backbone_0i_25_15 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[7]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[7]),.ZN(mem_backbone_0_n_25_8));
	INV_X1_LVT mem_backbone_0i_25_16 (.A(mem_backbone_0_n_25_8),.ZN(dmem_din[7]));
	AOI22_X1_LVT mem_backbone_0i_24_13 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[6]),.B1(dbg_mem_en),.B2(dbg_mem_dout[6]),.ZN(mem_backbone_0_n_24_7));
	INV_X1_LVT mem_backbone_0i_24_14 (.A(mem_backbone_0_n_24_7),.ZN(pmem_din[6]));
	AOI22_X1_LVT mem_backbone_0i_25_13 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[6]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[6]),.ZN(mem_backbone_0_n_25_7));
	INV_X1_LVT mem_backbone_0i_25_14 (.A(mem_backbone_0_n_25_7),.ZN(dmem_din[6]));
	AOI22_X1_LVT mem_backbone_0i_24_11 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[5]),.B1(dbg_mem_en),.B2(dbg_mem_dout[5]),.ZN(mem_backbone_0_n_24_6));
	INV_X1_LVT mem_backbone_0i_24_12 (.A(mem_backbone_0_n_24_6),.ZN(pmem_din[5]));
	AOI22_X1_LVT mem_backbone_0i_25_11 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[5]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[5]),.ZN(mem_backbone_0_n_25_6));
	INV_X1_LVT mem_backbone_0i_25_12 (.A(mem_backbone_0_n_25_6),.ZN(dmem_din[5]));
	AOI22_X1_LVT mem_backbone_0i_24_9 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[4]),.B1(dbg_mem_en),.B2(dbg_mem_dout[4]),.ZN(mem_backbone_0_n_24_5));
	INV_X1_LVT mem_backbone_0i_24_10 (.A(mem_backbone_0_n_24_5),.ZN(pmem_din[4]));
	AOI22_X1_LVT mem_backbone_0i_25_9 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[4]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[4]),.ZN(mem_backbone_0_n_25_5));
	INV_X1_LVT mem_backbone_0i_25_10 (.A(mem_backbone_0_n_25_5),.ZN(dmem_din[4]));
	AOI22_X1_LVT mem_backbone_0i_24_7 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[3]),.B1(dbg_mem_en),.B2(dbg_mem_dout[3]),.ZN(mem_backbone_0_n_24_4));
	INV_X1_LVT mem_backbone_0i_24_8 (.A(mem_backbone_0_n_24_4),.ZN(pmem_din[3]));
	AOI22_X1_LVT mem_backbone_0i_25_7 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[3]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[3]),.ZN(mem_backbone_0_n_25_4));
	INV_X1_LVT mem_backbone_0i_25_8 (.A(mem_backbone_0_n_25_4),.ZN(dmem_din[3]));
	AOI22_X1_LVT mem_backbone_0i_24_5 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[2]),.B1(dbg_mem_en),.B2(dbg_mem_dout[2]),.ZN(mem_backbone_0_n_24_3));
	INV_X1_LVT mem_backbone_0i_24_6 (.A(mem_backbone_0_n_24_3),.ZN(pmem_din[2]));
	AOI22_X1_LVT mem_backbone_0i_25_5 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[2]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[2]),.ZN(mem_backbone_0_n_25_3));
	INV_X1_LVT mem_backbone_0i_25_6 (.A(mem_backbone_0_n_25_3),.ZN(dmem_din[2]));
	AOI22_X1_LVT mem_backbone_0i_24_3 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[1]),.B1(dbg_mem_en),.B2(dbg_mem_dout[1]),.ZN(mem_backbone_0_n_24_2));
	INV_X1_LVT mem_backbone_0i_24_4 (.A(mem_backbone_0_n_24_2),.ZN(pmem_din[1]));
	AOI22_X1_LVT mem_backbone_0i_25_3 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[1]),.B1(mem_backbone_0_ext_dmem_en),.B2(pmem_din[1]),.ZN(mem_backbone_0_n_25_2));
	INV_X1_LVT mem_backbone_0i_25_4 (.A(mem_backbone_0_n_25_2),.ZN(dmem_din[1]));
	AOI22_X1_LVT mem_backbone_0i_24_1 (.A1(mem_backbone_0_n_24_0),.A2(dma_din[0]),.B1(dbg_mem_dout[0]),.B2(dbg_mem_en),.ZN(mem_backbone_0_n_24_1));
	INV_X1_LVT mem_backbone_0i_24_2 (.A(mem_backbone_0_n_24_1),.ZN(pmem_din[0]));
	AOI22_X1_LVT mem_backbone_0i_25_1 (.A1(mem_backbone_0_n_25_0),.A2(eu_mdb_out[0]),.B1(pmem_din[0]),.B2(mem_backbone_0_ext_dmem_en),.ZN(mem_backbone_0_n_25_1));
	INV_X1_LVT mem_backbone_0i_25_2 (.A(mem_backbone_0_n_25_1),.ZN(dmem_din[0]));
	INV_X1_LVT mem_backbone_0i_29_0 (.A(mem_backbone_0_ext_dmem_en),.ZN(mem_backbone_0_n_29_0));
	INV_X1_LVT mem_backbone_0i_26_1 (.A(eu_mb_wr[1]),.ZN(mem_backbone_0_n_8));
	INV_X1_LVT mem_backbone_0i_27_0 (.A(dbg_mem_en),.ZN(mem_backbone_0_n_27_0));
	AOI22_X1_LVT mem_backbone_0i_27_3 (.A1(mem_backbone_0_n_27_0),.A2(dma_we[1]),.B1(dbg_mem_en),.B2(dbg_mem_wr[1]),.ZN(mem_backbone_0_n_27_2));
	INV_X1_LVT mem_backbone_0i_27_4 (.A(mem_backbone_0_n_27_2),.ZN(mem_backbone_0_ext_mem_wr[1]));
	INV_X1_LVT mem_backbone_0i_28_1 (.A(mem_backbone_0_ext_mem_wr[1]),.ZN(mem_backbone_0_n_10));
	AOI22_X1_LVT mem_backbone_0i_29_3 (.A1(mem_backbone_0_n_29_0),.A2(mem_backbone_0_n_8),.B1(mem_backbone_0_ext_dmem_en),.B2(mem_backbone_0_n_10),.ZN(mem_backbone_0_n_29_2));
	INV_X1_LVT mem_backbone_0i_29_4 (.A(mem_backbone_0_n_29_2),.ZN(dmem_wen[1]));
	INV_X1_LVT mem_backbone_0i_26_0 (.A(eu_mb_wr[0]),.ZN(mem_backbone_0_n_7));
	AOI22_X1_LVT mem_backbone_0i_27_1 (.A1(mem_backbone_0_n_27_0),.A2(dma_we[0]),.B1(dbg_mem_wr[0]),.B2(dbg_mem_en),.ZN(mem_backbone_0_n_27_1));
	INV_X1_LVT mem_backbone_0i_27_2 (.A(mem_backbone_0_n_27_1),.ZN(mem_backbone_0_ext_mem_wr[0]));
	INV_X1_LVT mem_backbone_0i_28_0 (.A(mem_backbone_0_ext_mem_wr[0]),.ZN(mem_backbone_0_n_9));
	AOI22_X1_LVT mem_backbone_0i_29_1 (.A1(mem_backbone_0_n_29_0),.A2(mem_backbone_0_n_7),.B1(mem_backbone_0_n_9),.B2(mem_backbone_0_ext_dmem_en),.ZN(mem_backbone_0_n_29_1));
	INV_X1_LVT mem_backbone_0i_29_2 (.A(mem_backbone_0_n_29_1),.ZN(dmem_wen[0]));
	DFFR_X1_LVT mem_backbone_0eu_mdb_in_sel_reg___05F05b1___05F05d (.D(mem_backbone_0_eu_pmem_en),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_eu_mdb_in_sel[1]),.QN());
	DFFR_X1_LVT mem_backbone_0eu_mdb_in_sel_reg___05F05b0___05F05d (.D(mem_backbone_0_eu_per_en),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_eu_mdb_in_sel[0]),.QN());
	INV_X1_LVT mem_backbone_0i_31_1 (.A(mem_backbone_0_eu_mdb_in_sel[0]),.ZN(mem_backbone_0_n_31_0));
	NOR2_X1_LVT mem_backbone_0i_31_2 (.A1(mem_backbone_0_n_31_0),.A2(mem_backbone_0_eu_mdb_in_sel[1]),.ZN(mem_backbone_0_n_12));
	NOR2_X1_LVT mem_backbone_0i_31_0 (.A1(mem_backbone_0_eu_mdb_in_sel[0]),.A2(mem_backbone_0_eu_mdb_in_sel[1]),.ZN(mem_backbone_0_n_11));
	AOI222_X1_LVT mem_backbone_0i_32_30 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[15]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[15]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[15]),.ZN(mem_backbone_0_n_32_15));
	INV_X1_LVT mem_backbone_0i_32_31 (.A(mem_backbone_0_n_32_15),.ZN(eu_mdb_in[15]));
	AOI222_X1_LVT mem_backbone_0i_32_28 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[14]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[14]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[14]),.ZN(mem_backbone_0_n_32_14));
	INV_X1_LVT mem_backbone_0i_32_29 (.A(mem_backbone_0_n_32_14),.ZN(eu_mdb_in[14]));
	AOI222_X1_LVT mem_backbone_0i_32_26 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[13]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[13]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[13]),.ZN(mem_backbone_0_n_32_13));
	INV_X1_LVT mem_backbone_0i_32_27 (.A(mem_backbone_0_n_32_13),.ZN(eu_mdb_in[13]));
	AOI222_X1_LVT mem_backbone_0i_32_24 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[12]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[12]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[12]),.ZN(mem_backbone_0_n_32_12));
	INV_X1_LVT mem_backbone_0i_32_25 (.A(mem_backbone_0_n_32_12),.ZN(eu_mdb_in[12]));
	AOI222_X1_LVT mem_backbone_0i_32_22 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[11]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[11]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[11]),.ZN(mem_backbone_0_n_32_11));
	INV_X1_LVT mem_backbone_0i_32_23 (.A(mem_backbone_0_n_32_11),.ZN(eu_mdb_in[11]));
	AOI222_X1_LVT mem_backbone_0i_32_20 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[10]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[10]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[10]),.ZN(mem_backbone_0_n_32_10));
	INV_X1_LVT mem_backbone_0i_32_21 (.A(mem_backbone_0_n_32_10),.ZN(eu_mdb_in[10]));
	AOI222_X1_LVT mem_backbone_0i_32_18 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[9]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[9]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[9]),.ZN(mem_backbone_0_n_32_9));
	INV_X1_LVT mem_backbone_0i_32_19 (.A(mem_backbone_0_n_32_9),.ZN(eu_mdb_in[9]));
	AOI222_X1_LVT mem_backbone_0i_32_16 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[8]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[8]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[8]),.ZN(mem_backbone_0_n_32_8));
	INV_X1_LVT mem_backbone_0i_32_17 (.A(mem_backbone_0_n_32_8),.ZN(eu_mdb_in[8]));
	AOI222_X1_LVT mem_backbone_0i_32_14 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[7]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[7]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[7]),.ZN(mem_backbone_0_n_32_7));
	INV_X1_LVT mem_backbone_0i_32_15 (.A(mem_backbone_0_n_32_7),.ZN(eu_mdb_in[7]));
	AOI222_X1_LVT mem_backbone_0i_32_12 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[6]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[6]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[6]),.ZN(mem_backbone_0_n_32_6));
	INV_X1_LVT mem_backbone_0i_32_13 (.A(mem_backbone_0_n_32_6),.ZN(eu_mdb_in[6]));
	AOI222_X1_LVT mem_backbone_0i_32_10 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[5]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[5]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[5]),.ZN(mem_backbone_0_n_32_5));
	INV_X1_LVT mem_backbone_0i_32_11 (.A(mem_backbone_0_n_32_5),.ZN(eu_mdb_in[5]));
	AOI222_X1_LVT mem_backbone_0i_32_8 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[4]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[4]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[4]),.ZN(mem_backbone_0_n_32_4));
	INV_X1_LVT mem_backbone_0i_32_9 (.A(mem_backbone_0_n_32_4),.ZN(eu_mdb_in[4]));
	AOI222_X1_LVT mem_backbone_0i_32_6 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[3]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[3]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[3]),.ZN(mem_backbone_0_n_32_3));
	INV_X1_LVT mem_backbone_0i_32_7 (.A(mem_backbone_0_n_32_3),.ZN(eu_mdb_in[3]));
	AOI222_X1_LVT mem_backbone_0i_32_4 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[2]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[2]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[2]),.ZN(mem_backbone_0_n_32_2));
	INV_X1_LVT mem_backbone_0i_32_5 (.A(mem_backbone_0_n_32_2),.ZN(eu_mdb_in[2]));
	AOI222_X1_LVT mem_backbone_0i_32_2 (.A1(mem_backbone_0_eu_mdb_in_sel[1]),.A2(pmem_dout[1]),.B1(mem_backbone_0_n_12),.B2(mem_backbone_0_per_dout_val[1]),.C1(mem_backbone_0_n_11),.C2(dmem_dout[1]),.ZN(mem_backbone_0_n_32_1));
	INV_X1_LVT mem_backbone_0i_32_3 (.A(mem_backbone_0_n_32_1),.ZN(eu_mdb_in[1]));
	AOI222_X1_LVT mem_backbone_0i_32_0 (.A1(pmem_dout[0]),.A2(mem_backbone_0_eu_mdb_in_sel[1]),.B1(mem_backbone_0_per_dout_val[0]),.B2(mem_backbone_0_n_12),.C1(dmem_dout[0]),.C2(mem_backbone_0_n_11),.ZN(mem_backbone_0_n_32_0));
	INV_X1_LVT mem_backbone_0i_32_1 (.A(mem_backbone_0_n_32_0),.ZN(eu_mdb_in[0]));
	DFFR_X1_LVT mem_backbone_0fe_pmem_en_dly_reg (.D(mem_backbone_0_fe_pmem_en),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_fe_pmem_en_dly),.QN());
	NAND2_X1_LVT mem_backbone_0i_33_0 (.A1(mem_backbone_0_n_0),.A2(mem_backbone_0_fe_pmem_en_dly),.ZN(mem_backbone_0_n_33_0));
	NOR2_X1_LVT mem_backbone_0i_33_1 (.A1(mem_backbone_0_n_33_0),.A2(cpu_halt_st),.ZN(mem_backbone_0_fe_pmem_save));
	INV_X1_LVT mem_backbone_0i_35_0 (.A(cpu_halt_st),.ZN(mem_backbone_0_n_35_0));
	INV_X1_LVT mem_backbone_0i_35_1 (.A(mem_backbone_0_fe_pmem_en),.ZN(mem_backbone_0_n_35_1));
	OAI21_X1_LVT mem_backbone_0i_35_2 (.A(mem_backbone_0_n_35_0),.B1(mem_backbone_0_n_35_1),.B2(mem_backbone_0_fe_pmem_en_dly),.ZN(mem_backbone_0_fe_pmem_restore));
	INV_X1_LVT mem_backbone_0i_37_1 (.A(mem_backbone_0_fe_pmem_restore),.ZN(mem_backbone_0_n_37_1));
	INV_X1_LVT mem_backbone_0i_37_0 (.A(mem_backbone_0_fe_pmem_save),.ZN(mem_backbone_0_n_37_0));
	NAND2_X1_LVT mem_backbone_0i_37_2 (.A1(mem_backbone_0_n_37_1),.A2(mem_backbone_0_n_37_0),.ZN(mem_backbone_0_n_15));
	CLKGATETST_X1_LVT mem_backbone_0clk_gate_pmem_dout_bckup_sel_reg (.CK(mclk),.E(mem_backbone_0_n_15),.SE(1'b0),.GCK(mem_backbone_0_n_14));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_sel_reg (.D(mem_backbone_0_fe_pmem_save),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_14),.Q(mem_backbone_0_pmem_dout_bckup_sel),.QN());
	INV_X1_LVT mem_backbone_0i_39_0 (.A(mem_backbone_0_pmem_dout_bckup_sel),.ZN(mem_backbone_0_n_39_0));
	CLKGATETST_X1_LVT mem_backbone_0clk_gate_pmem_dout_bckup_reg (.CK(mclk),.E(mem_backbone_0_fe_pmem_save),.SE(1'b0),.GCK(mem_backbone_0_n_13));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b15___05F05d (.D(pmem_dout[15]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[15]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_31 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[15]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[15]),.ZN(mem_backbone_0_n_39_16));
	INV_X1_LVT mem_backbone_0i_39_32 (.A(mem_backbone_0_n_39_16),.ZN(fe_mdb_in[15]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b14___05F05d (.D(pmem_dout[14]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[14]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_29 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[14]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[14]),.ZN(mem_backbone_0_n_39_15));
	INV_X1_LVT mem_backbone_0i_39_30 (.A(mem_backbone_0_n_39_15),.ZN(fe_mdb_in[14]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b13___05F05d (.D(pmem_dout[13]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[13]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_27 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[13]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[13]),.ZN(mem_backbone_0_n_39_14));
	INV_X1_LVT mem_backbone_0i_39_28 (.A(mem_backbone_0_n_39_14),.ZN(fe_mdb_in[13]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b12___05F05d (.D(pmem_dout[12]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[12]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_25 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[12]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[12]),.ZN(mem_backbone_0_n_39_13));
	INV_X1_LVT mem_backbone_0i_39_26 (.A(mem_backbone_0_n_39_13),.ZN(fe_mdb_in[12]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b11___05F05d (.D(pmem_dout[11]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[11]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_23 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[11]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[11]),.ZN(mem_backbone_0_n_39_12));
	INV_X1_LVT mem_backbone_0i_39_24 (.A(mem_backbone_0_n_39_12),.ZN(fe_mdb_in[11]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b10___05F05d (.D(pmem_dout[10]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[10]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_21 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[10]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[10]),.ZN(mem_backbone_0_n_39_11));
	INV_X1_LVT mem_backbone_0i_39_22 (.A(mem_backbone_0_n_39_11),.ZN(fe_mdb_in[10]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b9___05F05d (.D(pmem_dout[9]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[9]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_19 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[9]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[9]),.ZN(mem_backbone_0_n_39_10));
	INV_X1_LVT mem_backbone_0i_39_20 (.A(mem_backbone_0_n_39_10),.ZN(fe_mdb_in[9]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b8___05F05d (.D(pmem_dout[8]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[8]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_17 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[8]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[8]),.ZN(mem_backbone_0_n_39_9));
	INV_X1_LVT mem_backbone_0i_39_18 (.A(mem_backbone_0_n_39_9),.ZN(fe_mdb_in[8]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b7___05F05d (.D(pmem_dout[7]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[7]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_15 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[7]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[7]),.ZN(mem_backbone_0_n_39_8));
	INV_X1_LVT mem_backbone_0i_39_16 (.A(mem_backbone_0_n_39_8),.ZN(fe_mdb_in[7]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b6___05F05d (.D(pmem_dout[6]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[6]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_13 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[6]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[6]),.ZN(mem_backbone_0_n_39_7));
	INV_X1_LVT mem_backbone_0i_39_14 (.A(mem_backbone_0_n_39_7),.ZN(fe_mdb_in[6]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b5___05F05d (.D(pmem_dout[5]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[5]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_11 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[5]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[5]),.ZN(mem_backbone_0_n_39_6));
	INV_X1_LVT mem_backbone_0i_39_12 (.A(mem_backbone_0_n_39_6),.ZN(fe_mdb_in[5]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b4___05F05d (.D(pmem_dout[4]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[4]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_9 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[4]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[4]),.ZN(mem_backbone_0_n_39_5));
	INV_X1_LVT mem_backbone_0i_39_10 (.A(mem_backbone_0_n_39_5),.ZN(fe_mdb_in[4]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b3___05F05d (.D(pmem_dout[3]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[3]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_7 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[3]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[3]),.ZN(mem_backbone_0_n_39_4));
	INV_X1_LVT mem_backbone_0i_39_8 (.A(mem_backbone_0_n_39_4),.ZN(fe_mdb_in[3]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b2___05F05d (.D(pmem_dout[2]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[2]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_5 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[2]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[2]),.ZN(mem_backbone_0_n_39_3));
	INV_X1_LVT mem_backbone_0i_39_6 (.A(mem_backbone_0_n_39_3),.ZN(fe_mdb_in[2]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b1___05F05d (.D(pmem_dout[1]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[1]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_3 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[1]),.B1(mem_backbone_0_pmem_dout_bckup_sel),.B2(mem_backbone_0_pmem_dout_bckup[1]),.ZN(mem_backbone_0_n_39_2));
	INV_X1_LVT mem_backbone_0i_39_4 (.A(mem_backbone_0_n_39_2),.ZN(fe_mdb_in[1]));
	DFFR_X1_LVT mem_backbone_0pmem_dout_bckup_reg___05F05b0___05F05d (.D(pmem_dout[0]),.RN(mem_backbone_0_n_2),.CK(mem_backbone_0_n_13),.Q(mem_backbone_0_pmem_dout_bckup[0]),.QN());
	AOI22_X1_LVT mem_backbone_0i_39_1 (.A1(mem_backbone_0_n_39_0),.A2(pmem_dout[0]),.B1(mem_backbone_0_pmem_dout_bckup[0]),.B2(mem_backbone_0_pmem_dout_bckup_sel),.ZN(mem_backbone_0_n_39_1));
	INV_X1_LVT mem_backbone_0i_39_2 (.A(mem_backbone_0_n_39_1),.ZN(fe_mdb_in[0]));
	AND2_X1_LVT mem_backbone_0i_40_0 (.A1(mem_backbone_0_fe_pmem_en),.A2(mem_backbone_0_eu_pmem_en),.ZN(fe_pmem_wait));
	INV_X1_LVT mem_backbone_0i_41_0 (.A(dbg_mem_en),.ZN(mem_backbone_0_n_16));
	NAND2_X1_LVT mem_backbone_0i_42_0 (.A1(mem_backbone_0_n_16),.A2(dma_en),.ZN(mem_backbone_0_n_42_0));
	NOR4_X1_LVT mem_backbone_0i_42_1 (.A1(mem_backbone_0_n_42_0),.A2(mem_backbone_0_ext_dmem_sel),.A3(mem_backbone_0_ext_per_sel),.A4(mem_backbone_0_ext_pmem_sel),.ZN(dma_resp));
	OR4_X1_LVT mem_backbone_0i_43_0 (.A1(mem_backbone_0_ext_dmem_en),.A2(dma_resp),.A3(mem_backbone_0_ext_per_en),.A4(mem_backbone_0_ext_pmem_en),.ZN(mem_backbone_0_n_43_0));
	AND2_X1_LVT mem_backbone_0i_43_1 (.A1(mem_backbone_0_n_43_0),.A2(mem_backbone_0_n_16),.ZN(dma_ready));
	DFFR_X1_LVT mem_backbone_0dma_ready_dly_reg (.D(dma_ready),.RN(mem_backbone_0_n_2),.CK(mclk),.Q(mem_backbone_0_dma_ready_dly),.QN());
	AND2_X1_LVT mem_backbone_0i_44_15 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[15]),.ZN(dma_dout[15]));
	AND2_X1_LVT mem_backbone_0i_44_14 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[14]),.ZN(dma_dout[14]));
	AND2_X1_LVT mem_backbone_0i_44_13 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[13]),.ZN(dma_dout[13]));
	AND2_X1_LVT mem_backbone_0i_44_12 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[12]),.ZN(dma_dout[12]));
	AND2_X1_LVT mem_backbone_0i_44_11 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[11]),.ZN(dma_dout[11]));
	AND2_X1_LVT mem_backbone_0i_44_10 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[10]),.ZN(dma_dout[10]));
	AND2_X1_LVT mem_backbone_0i_44_9 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[9]),.ZN(dma_dout[9]));
	AND2_X1_LVT mem_backbone_0i_44_8 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[8]),.ZN(dma_dout[8]));
	AND2_X1_LVT mem_backbone_0i_44_7 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[7]),.ZN(dma_dout[7]));
	AND2_X1_LVT mem_backbone_0i_44_6 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[6]),.ZN(dma_dout[6]));
	AND2_X1_LVT mem_backbone_0i_44_5 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[5]),.ZN(dma_dout[5]));
	AND2_X1_LVT mem_backbone_0i_44_4 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[4]),.ZN(dma_dout[4]));
	AND2_X1_LVT mem_backbone_0i_44_3 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[3]),.ZN(dma_dout[3]));
	AND2_X1_LVT mem_backbone_0i_44_2 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[2]),.ZN(dma_dout[2]));
	AND2_X1_LVT mem_backbone_0i_44_1 (.A1(mem_backbone_0_dma_ready_dly),.A2(dbg_mem_din[1]),.ZN(dma_dout[1]));
	AND2_X1_LVT mem_backbone_0i_44_0 (.A1(dbg_mem_din[0]),.A2(mem_backbone_0_dma_ready_dly),.ZN(dma_dout[0]));
	INV_X1_LVT mem_backbone_0i_45_0 (.A(mem_backbone_0_ext_per_en),.ZN(mem_backbone_0_n_45_0));
	AOI22_X1_LVT mem_backbone_0i_45_15 (.A1(mem_backbone_0_n_45_0),.A2(eu_mab[8]),.B1(mem_backbone_0_ext_per_en),.B2(mem_backbone_0_ext_mem_addr[7]),.ZN(mem_backbone_0_n_45_8));
	INV_X1_LVT mem_backbone_0i_45_16 (.A(mem_backbone_0_n_45_8),.ZN(per_addr[7]));
	AOI22_X1_LVT mem_backbone_0i_45_13 (.A1(mem_backbone_0_n_45_0),.A2(eu_mab[7]),.B1(mem_backbone_0_ext_per_en),.B2(mem_backbone_0_ext_mem_addr[6]),.ZN(mem_backbone_0_n_45_7));
	INV_X1_LVT mem_backbone_0i_45_14 (.A(mem_backbone_0_n_45_7),.ZN(per_addr[6]));
	AOI22_X1_LVT mem_backbone_0i_45_11 (.A1(mem_backbone_0_n_45_0),.A2(eu_mab[6]),.B1(mem_backbone_0_ext_per_en),.B2(mem_backbone_0_ext_mem_addr[5]),.ZN(mem_backbone_0_n_45_6));
	INV_X1_LVT mem_backbone_0i_45_12 (.A(mem_backbone_0_n_45_6),.ZN(per_addr[5]));
	AOI22_X1_LVT mem_backbone_0i_45_9 (.A1(mem_backbone_0_n_45_0),.A2(eu_mab[5]),.B1(mem_backbone_0_ext_per_en),.B2(mem_backbone_0_ext_mem_addr[4]),.ZN(mem_backbone_0_n_45_5));
	INV_X1_LVT mem_backbone_0i_45_10 (.A(mem_backbone_0_n_45_5),.ZN(per_addr[4]));
	AOI22_X1_LVT mem_backbone_0i_45_7 (.A1(mem_backbone_0_n_45_0),.A2(eu_mab[4]),.B1(mem_backbone_0_ext_per_en),.B2(mem_backbone_0_ext_mem_addr[3]),.ZN(mem_backbone_0_n_45_4));
	INV_X1_LVT mem_backbone_0i_45_8 (.A(mem_backbone_0_n_45_4),.ZN(per_addr[3]));
	AOI22_X1_LVT mem_backbone_0i_45_5 (.A1(mem_backbone_0_n_45_0),.A2(eu_mab[3]),.B1(mem_backbone_0_ext_per_en),.B2(mem_backbone_0_ext_mem_addr[2]),.ZN(mem_backbone_0_n_45_3));
	INV_X1_LVT mem_backbone_0i_45_6 (.A(mem_backbone_0_n_45_3),.ZN(per_addr[2]));
	AOI22_X1_LVT mem_backbone_0i_45_3 (.A1(mem_backbone_0_n_45_0),.A2(eu_mab[2]),.B1(mem_backbone_0_ext_per_en),.B2(mem_backbone_0_ext_mem_addr[1]),.ZN(mem_backbone_0_n_45_2));
	INV_X1_LVT mem_backbone_0i_45_4 (.A(mem_backbone_0_n_45_2),.ZN(per_addr[1]));
	AOI22_X1_LVT mem_backbone_0i_45_1 (.A1(mem_backbone_0_n_45_0),.A2(eu_mab[1]),.B1(mem_backbone_0_ext_mem_addr[0]),.B2(mem_backbone_0_ext_per_en),.ZN(mem_backbone_0_n_45_1));
	INV_X1_LVT mem_backbone_0i_45_2 (.A(mem_backbone_0_n_45_1),.ZN(per_addr[0]));
	INV_X1_LVT mem_backbone_0i_46_0 (.A(mem_backbone_0_ext_per_en),.ZN(mem_backbone_0_n_46_0));
	AOI22_X1_LVT mem_backbone_0i_46_31 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[15]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[15]),.ZN(mem_backbone_0_n_46_16));
	INV_X1_LVT mem_backbone_0i_46_32 (.A(mem_backbone_0_n_46_16),.ZN(per_din[15]));
	AOI22_X1_LVT mem_backbone_0i_46_29 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[14]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[14]),.ZN(mem_backbone_0_n_46_15));
	INV_X1_LVT mem_backbone_0i_46_30 (.A(mem_backbone_0_n_46_15),.ZN(per_din[14]));
	AOI22_X1_LVT mem_backbone_0i_46_27 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[13]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[13]),.ZN(mem_backbone_0_n_46_14));
	INV_X1_LVT mem_backbone_0i_46_28 (.A(mem_backbone_0_n_46_14),.ZN(per_din[13]));
	AOI22_X1_LVT mem_backbone_0i_46_25 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[12]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[12]),.ZN(mem_backbone_0_n_46_13));
	INV_X1_LVT mem_backbone_0i_46_26 (.A(mem_backbone_0_n_46_13),.ZN(per_din[12]));
	AOI22_X1_LVT mem_backbone_0i_46_23 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[11]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[11]),.ZN(mem_backbone_0_n_46_12));
	INV_X1_LVT mem_backbone_0i_46_24 (.A(mem_backbone_0_n_46_12),.ZN(per_din[11]));
	AOI22_X1_LVT mem_backbone_0i_46_21 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[10]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[10]),.ZN(mem_backbone_0_n_46_11));
	INV_X1_LVT mem_backbone_0i_46_22 (.A(mem_backbone_0_n_46_11),.ZN(per_din[10]));
	AOI22_X1_LVT mem_backbone_0i_46_19 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[9]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[9]),.ZN(mem_backbone_0_n_46_10));
	INV_X1_LVT mem_backbone_0i_46_20 (.A(mem_backbone_0_n_46_10),.ZN(per_din[9]));
	AOI22_X1_LVT mem_backbone_0i_46_17 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[8]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[8]),.ZN(mem_backbone_0_n_46_9));
	INV_X1_LVT mem_backbone_0i_46_18 (.A(mem_backbone_0_n_46_9),.ZN(per_din[8]));
	AOI22_X1_LVT mem_backbone_0i_46_15 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[7]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[7]),.ZN(mem_backbone_0_n_46_8));
	INV_X1_LVT mem_backbone_0i_46_16 (.A(mem_backbone_0_n_46_8),.ZN(per_din[7]));
	AOI22_X1_LVT mem_backbone_0i_46_13 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[6]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[6]),.ZN(mem_backbone_0_n_46_7));
	INV_X1_LVT mem_backbone_0i_46_14 (.A(mem_backbone_0_n_46_7),.ZN(per_din[6]));
	AOI22_X1_LVT mem_backbone_0i_46_11 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[5]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[5]),.ZN(mem_backbone_0_n_46_6));
	INV_X1_LVT mem_backbone_0i_46_12 (.A(mem_backbone_0_n_46_6),.ZN(per_din[5]));
	AOI22_X1_LVT mem_backbone_0i_46_9 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[4]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[4]),.ZN(mem_backbone_0_n_46_5));
	INV_X1_LVT mem_backbone_0i_46_10 (.A(mem_backbone_0_n_46_5),.ZN(per_din[4]));
	AOI22_X1_LVT mem_backbone_0i_46_7 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[3]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[3]),.ZN(mem_backbone_0_n_46_4));
	INV_X1_LVT mem_backbone_0i_46_8 (.A(mem_backbone_0_n_46_4),.ZN(per_din[3]));
	AOI22_X1_LVT mem_backbone_0i_46_5 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[2]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[2]),.ZN(mem_backbone_0_n_46_3));
	INV_X1_LVT mem_backbone_0i_46_6 (.A(mem_backbone_0_n_46_3),.ZN(per_din[2]));
	AOI22_X1_LVT mem_backbone_0i_46_3 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[1]),.B1(mem_backbone_0_ext_per_en),.B2(pmem_din[1]),.ZN(mem_backbone_0_n_46_2));
	INV_X1_LVT mem_backbone_0i_46_4 (.A(mem_backbone_0_n_46_2),.ZN(per_din[1]));
	AOI22_X1_LVT mem_backbone_0i_46_1 (.A1(mem_backbone_0_n_46_0),.A2(eu_mdb_out[0]),.B1(pmem_din[0]),.B2(mem_backbone_0_ext_per_en),.ZN(mem_backbone_0_n_46_1));
	INV_X1_LVT mem_backbone_0i_46_2 (.A(mem_backbone_0_n_46_1),.ZN(per_din[0]));
	INV_X1_LVT mem_backbone_0i_47_0 (.A(mem_backbone_0_ext_per_en),.ZN(mem_backbone_0_n_47_0));
	AOI22_X1_LVT mem_backbone_0i_47_3 (.A1(mem_backbone_0_n_47_0),.A2(eu_mb_wr[1]),.B1(mem_backbone_0_ext_per_en),.B2(mem_backbone_0_ext_mem_wr[1]),.ZN(mem_backbone_0_n_47_2));
	INV_X1_LVT mem_backbone_0i_47_4 (.A(mem_backbone_0_n_47_2),.ZN(per_we[1]));
	AOI22_X1_LVT mem_backbone_0i_47_1 (.A1(mem_backbone_0_n_47_0),.A2(eu_mb_wr[0]),.B1(mem_backbone_0_ext_mem_wr[0]),.B2(mem_backbone_0_ext_per_en),.ZN(mem_backbone_0_n_47_1));
	INV_X1_LVT mem_backbone_0i_47_2 (.A(mem_backbone_0_n_47_1),.ZN(per_we[0]));
	OR2_X1_LVT mem_backbone_0i_48_0 (.A1(mem_backbone_0_ext_per_en),.A2(mem_backbone_0_eu_per_en),.ZN(per_en));
	NOR2_X1_LVT mem_backbone_0i_49_0 (.A1(mem_backbone_0_eu_pmem_en),.A2(mem_backbone_0_ext_pmem_en),.ZN(mem_backbone_0_n_49_0));
	AOI222_X1_LVT mem_backbone_0i_49_21 (.A1(mem_backbone_0_n_49_0),.A2(n_4),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[10]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[11]),.ZN(mem_backbone_0_n_49_11));
	INV_X1_LVT mem_backbone_0i_49_22 (.A(mem_backbone_0_n_49_11),.ZN(pmem_addr[10]));
	AOI222_X1_LVT mem_backbone_0i_49_19 (.A1(mem_backbone_0_n_49_0),.A2(n_5),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[9]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[10]),.ZN(mem_backbone_0_n_49_10));
	INV_X1_LVT mem_backbone_0i_49_20 (.A(mem_backbone_0_n_49_10),.ZN(pmem_addr[9]));
	AOI222_X1_LVT mem_backbone_0i_49_17 (.A1(mem_backbone_0_n_49_0),.A2(n_6),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[8]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[9]),.ZN(mem_backbone_0_n_49_9));
	INV_X1_LVT mem_backbone_0i_49_18 (.A(mem_backbone_0_n_49_9),.ZN(pmem_addr[8]));
	AOI222_X1_LVT mem_backbone_0i_49_15 (.A1(mem_backbone_0_n_49_0),.A2(n_7),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[7]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[8]),.ZN(mem_backbone_0_n_49_8));
	INV_X1_LVT mem_backbone_0i_49_16 (.A(mem_backbone_0_n_49_8),.ZN(pmem_addr[7]));
	AOI222_X1_LVT mem_backbone_0i_49_13 (.A1(mem_backbone_0_n_49_0),.A2(n_8),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[6]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[7]),.ZN(mem_backbone_0_n_49_7));
	INV_X1_LVT mem_backbone_0i_49_14 (.A(mem_backbone_0_n_49_7),.ZN(pmem_addr[6]));
	AOI222_X1_LVT mem_backbone_0i_49_11 (.A1(mem_backbone_0_n_49_0),.A2(n_9),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[5]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[6]),.ZN(mem_backbone_0_n_49_6));
	INV_X1_LVT mem_backbone_0i_49_12 (.A(mem_backbone_0_n_49_6),.ZN(pmem_addr[5]));
	AOI222_X1_LVT mem_backbone_0i_49_9 (.A1(mem_backbone_0_n_49_0),.A2(n_10),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[4]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[5]),.ZN(mem_backbone_0_n_49_5));
	INV_X1_LVT mem_backbone_0i_49_10 (.A(mem_backbone_0_n_49_5),.ZN(pmem_addr[4]));
	AOI222_X1_LVT mem_backbone_0i_49_7 (.A1(mem_backbone_0_n_49_0),.A2(n_11),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[3]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[4]),.ZN(mem_backbone_0_n_49_4));
	INV_X1_LVT mem_backbone_0i_49_8 (.A(mem_backbone_0_n_49_4),.ZN(pmem_addr[3]));
	AOI222_X1_LVT mem_backbone_0i_49_5 (.A1(mem_backbone_0_n_49_0),.A2(n_12),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[2]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[3]),.ZN(mem_backbone_0_n_49_3));
	INV_X1_LVT mem_backbone_0i_49_6 (.A(mem_backbone_0_n_49_3),.ZN(pmem_addr[2]));
	AOI222_X1_LVT mem_backbone_0i_49_3 (.A1(mem_backbone_0_n_49_0),.A2(n_13),.B1(mem_backbone_0_ext_pmem_en),.B2(mem_backbone_0_ext_mem_addr[1]),.C1(mem_backbone_0_eu_pmem_en),.C2(eu_mab[2]),.ZN(mem_backbone_0_n_49_2));
	INV_X1_LVT mem_backbone_0i_49_4 (.A(mem_backbone_0_n_49_2),.ZN(pmem_addr[1]));
	AOI222_X1_LVT mem_backbone_0i_49_1 (.A1(mem_backbone_0_n_49_0),.A2(n_14),.B1(mem_backbone_0_ext_mem_addr[0]),.B2(mem_backbone_0_ext_pmem_en),.C1(eu_mab[1]),.C2(mem_backbone_0_eu_pmem_en),.ZN(mem_backbone_0_n_49_1));
	INV_X1_LVT mem_backbone_0i_49_2 (.A(mem_backbone_0_n_49_1),.ZN(pmem_addr[0]));
	NOR3_X1_LVT mem_backbone_0i_50_0 (.A1(mem_backbone_0_fe_pmem_en),.A2(mem_backbone_0_ext_pmem_en),.A3(mem_backbone_0_eu_pmem_en),.ZN(pmem_cen));
	NAND2_X1_LVT mem_backbone_0i_51_2 (.A1(mem_backbone_0_ext_pmem_en),.A2(mem_backbone_0_n_10),.ZN(mem_backbone_0_n_51_1));
	NAND2_X1_LVT mem_backbone_0i_51_3 (.A1(mem_backbone_0_n_51_1),.A2(mem_backbone_0_ext_pmem_en),.ZN(pmem_wen[1]));
	NAND2_X1_LVT mem_backbone_0i_51_0 (.A1(mem_backbone_0_n_9),.A2(mem_backbone_0_ext_pmem_en),.ZN(mem_backbone_0_n_51_0));
	NAND2_X1_LVT mem_backbone_0i_51_1 (.A1(mem_backbone_0_n_51_0),.A2(mem_backbone_0_ext_pmem_en),.ZN(pmem_wen[0]));
	INV_X1_LVT frontend_0i_78_0 (.A(puc_rst),.ZN(frontend_0_n_91));
	DFFR_X1_LVT frontend_0i_state_reg___05F05b0___05F05d (.D(frontend_0_i_state_nxt_reg[0]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(frontend_0_i_state[0]),.QN());
	INV_X1_LVT frontend_0i_76_2 (.A(frontend_0_i_state[0]),.ZN(frontend_0_n_76_2));
	INV_X1_LVT frontend_0i_76_1 (.A(frontend_0_i_state[2]),.ZN(frontend_0_n_76_1));
	NOR3_X1_LVT frontend_0i_76_3 (.A1(frontend_0_n_76_1),.A2(frontend_0_n_76_2),.A3(frontend_0_i_state[1]),.ZN(frontend_0_n_76_3));
	INV_X1_LVT frontend_0i_0_0 (.A(cpu_halt_cmd),.ZN(frontend_0_n_0_0));
	NAND2_X1_LVT frontend_0i_0_1 (.A1(frontend_0_n_0_0),.A2(cpu_en_s),.ZN(frontend_0_cpu_halt_req));
	INV_X1_LVT frontend_0i_1_0 (.A(frontend_0_cpu_halt_req),.ZN(frontend_0_n_0));
	INV_X1_LVT frontend_0i_74_0 (.A(frontend_0_n_0),.ZN(frontend_0_n_74_0));
	NOR2_X1_LVT frontend_0i_74_1 (.A1(frontend_0_n_74_0),.A2(cpuoff),.ZN(frontend_0_n_87));
	INV_X1_LVT frontend_0i_2_0 (.A(cpu_halt_st),.ZN(frontend_0_n_1));
	NAND2_X1_LVT frontend_0i_4_0 (.A1(frontend_0_n_1),.A2(frontend_0_n_0),.ZN(frontend_0_n_4_0));
	NOR4_X1_LVT frontend_0i_3_0 (.A1(irq[10]),.A2(irq[11]),.A3(irq[12]),.A4(irq[13]),.ZN(frontend_0_n_3_0));
	NOR4_X1_LVT frontend_0i_3_1 (.A1(irq[2]),.A2(irq[3]),.A3(irq[4]),.A4(irq[5]),.ZN(frontend_0_n_3_1));
	NOR4_X1_LVT frontend_0i_3_2 (.A1(irq[6]),.A2(irq[7]),.A3(irq[8]),.A4(irq[9]),.ZN(frontend_0_n_3_2));
	NOR2_X1_LVT frontend_0i_3_3 (.A1(irq[0]),.A2(irq[1]),.ZN(frontend_0_n_3_3));
	NAND4_X1_LVT frontend_0i_3_4 (.A1(frontend_0_n_3_0),.A2(frontend_0_n_3_1),.A3(frontend_0_n_3_2),.A4(frontend_0_n_3_3),.ZN(frontend_0_n_2));
	OAI21_X1_LVT frontend_0i_4_1 (.A(gie),.B1(frontend_0_n_2),.B2(wdt_irq),.ZN(frontend_0_n_4_1));
	INV_X1_LVT frontend_0i_4_2 (.A(nmi_pnd),.ZN(frontend_0_n_4_2));
	AOI21_X1_LVT frontend_0i_4_3 (.A(frontend_0_n_4_0),.B1(frontend_0_n_4_1),.B2(frontend_0_n_4_2),.ZN(frontend_0_n_3));
	AND2_X1_LVT frontend_0i_74_2 (.A1(frontend_0_n_0),.A2(frontend_0_n_3),.ZN(frontend_0_n_88));
	NOR2_X1_LVT frontend_0i_75_0 (.A1(frontend_0_n_87),.A2(frontend_0_n_88),.ZN(frontend_0_n_89));
	AND2_X1_LVT frontend_0i_76_4 (.A1(frontend_0_n_76_3),.A2(frontend_0_n_89),.ZN(frontend_0_n_76_4));
	INV_X1_LVT frontend_0i_76_5 (.A(frontend_0_i_state[1]),.ZN(frontend_0_n_76_5));
	NOR3_X1_LVT frontend_0i_76_6 (.A1(frontend_0_n_76_5),.A2(frontend_0_i_state[0]),.A3(frontend_0_i_state[2]),.ZN(frontend_0_n_76_6));
	INV_X1_LVT frontend_0i_55_0 (.A(e_state[0]),.ZN(frontend_0_n_55_0));
	INV_X1_LVT frontend_0i_6_2 (.A(frontend_0_i_state[2]),.ZN(frontend_0_n_6_1));
	INV_X1_LVT frontend_0i_6_3 (.A(frontend_0_i_state[0]),.ZN(frontend_0_n_6_2));
	NOR3_X1_LVT frontend_0i_6_4 (.A1(frontend_0_n_6_1),.A2(frontend_0_n_6_2),.A3(frontend_0_i_state[1]),.ZN(frontend_0_n_5));
	OR2_X1_LVT frontend_0i_49_2 (.A1(frontend_0_n_5),.A2(frontend_0_cpu_halt_req),.ZN(frontend_0_n_55));
	NOR3_X1_LVT frontend_0i_8_0 (.A1(fe_mdb_in[13]),.A2(fe_mdb_in[14]),.A3(fe_mdb_in[15]),.ZN(frontend_0_n_10));
	NAND2_X1_LVT frontend_0i_25_5 (.A1(fe_mdb_in[7]),.A2(fe_mdb_in[8]),.ZN(frontend_0_n_25_5));
	INV_X1_LVT frontend_0i_25_6 (.A(fe_mdb_in[9]),.ZN(frontend_0_n_25_6));
	NOR2_X1_LVT frontend_0i_25_14 (.A1(frontend_0_n_25_5),.A2(frontend_0_n_25_6),.ZN(frontend_0_n_29));
	AND2_X1_LVT frontend_0i_26_7 (.A1(frontend_0_n_10),.A2(frontend_0_n_29),.ZN(frontend_0_n_37));
	INV_X1_LVT frontend_0i_27_8 (.A(frontend_0_n_37),.ZN(frontend_0_n_27_1));
	INV_X1_LVT frontend_0i_25_0 (.A(fe_mdb_in[7]),.ZN(frontend_0_n_25_0));
	NAND2_X1_LVT frontend_0i_25_4 (.A1(frontend_0_n_25_0),.A2(fe_mdb_in[8]),.ZN(frontend_0_n_25_4));
	NOR2_X1_LVT frontend_0i_25_13 (.A1(frontend_0_n_25_4),.A2(frontend_0_n_25_6),.ZN(frontend_0_n_28));
	AND2_X1_LVT frontend_0i_26_6 (.A1(frontend_0_n_10),.A2(frontend_0_n_28),.ZN(frontend_0_n_36));
	AND2_X1_LVT frontend_0i_27_7 (.A1(frontend_0_n_27_0),.A2(frontend_0_n_36),.ZN(frontend_0_inst_so_nxt[6]));
	INV_X1_LVT frontend_0i_7_0 (.A(frontend_0_irq_detect),.ZN(frontend_0_n_9));
	NAND2_X1_LVT frontend_0i_11_0 (.A1(fe_mdb_in[13]),.A2(frontend_0_n_9),.ZN(frontend_0_n_11_0));
	NOR3_X1_LVT frontend_0i_11_1 (.A1(frontend_0_n_11_0),.A2(fe_mdb_in[14]),.A3(fe_mdb_in[15]),.ZN(frontend_0_inst_type_nxt));
	OR2_X1_LVT frontend_0i_42_0 (.A1(frontend_0_inst_so_nxt[6]),.A2(frontend_0_inst_type_nxt),.ZN(frontend_0_n_49));
	INV_X1_LVT frontend_0i_23_0 (.A(fe_mdb_in[7]),.ZN(frontend_0_n_23_0));
	NOR4_X1_LVT frontend_0i_23_1 (.A1(frontend_0_n_23_0),.A2(fe_mdb_in[1]),.A3(fe_mdb_in[2]),.A4(fe_mdb_in[3]),.ZN(frontend_0_n_23_1));
	INV_X1_LVT frontend_0i_23_2 (.A(fe_mdb_in[0]),.ZN(frontend_0_n_23_2));
	NAND2_X1_LVT frontend_0i_23_3 (.A1(frontend_0_n_23_1),.A2(frontend_0_n_23_2),.ZN(frontend_0_n_23_3));
	NOR4_X1_LVT frontend_0i_23_4 (.A1(fe_mdb_in[0]),.A2(fe_mdb_in[1]),.A3(fe_mdb_in[2]),.A4(fe_mdb_in[3]),.ZN(frontend_0_n_23_4));
	INV_X1_LVT frontend_0i_23_5 (.A(frontend_0_n_23_4),.ZN(frontend_0_n_23_5));
	NAND2_X1_LVT frontend_0i_23_6 (.A1(frontend_0_n_23_3),.A2(frontend_0_n_23_5),.ZN(frontend_0_n_23_6));
	INV_X1_LVT frontend_0i_23_7 (.A(frontend_0_n_23_6),.ZN(frontend_0_n_23_7));
	AOI22_X1_LVT frontend_0i_23_8 (.A1(frontend_0_n_23_3),.A2(frontend_0_n_23_4),.B1(frontend_0_n_23_7),.B2(frontend_0_n_23_0),.ZN(frontend_0_n_23_8));
	INV_X1_LVT frontend_0i_23_9 (.A(fe_mdb_in[2]),.ZN(frontend_0_n_23_9));
	INV_X1_LVT frontend_0i_23_10 (.A(fe_mdb_in[3]),.ZN(frontend_0_n_23_10));
	NAND4_X1_LVT frontend_0i_23_11 (.A1(frontend_0_n_23_9),.A2(frontend_0_n_23_10),.A3(fe_mdb_in[7]),.A4(fe_mdb_in[1]),.ZN(frontend_0_n_23_11));
	OR2_X1_LVT frontend_0i_23_12 (.A1(frontend_0_n_23_11),.A2(fe_mdb_in[0]),.ZN(frontend_0_n_23_12));
	OAI21_X1_LVT frontend_0i_22_0 (.A(frontend_0_n_9),.B1(fe_mdb_in[14]),.B2(fe_mdb_in[15]),.ZN(frontend_0_n_22_0));
	INV_X1_LVT frontend_0i_22_1 (.A(frontend_0_n_22_0),.ZN(frontend_0_n_17));
	NAND2_X1_LVT frontend_0i_23_13 (.A1(frontend_0_n_23_12),.A2(frontend_0_n_17),.ZN(frontend_0_n_23_13));
	INV_X1_LVT frontend_0i_23_14 (.A(frontend_0_n_23_13),.ZN(frontend_0_n_23_14));
	NAND4_X1_LVT frontend_0i_23_15 (.A1(frontend_0_n_23_2),.A2(frontend_0_n_23_9),.A3(frontend_0_n_23_10),.A4(fe_mdb_in[1]),.ZN(frontend_0_n_23_15));
	NAND2_X1_LVT frontend_0i_23_16 (.A1(frontend_0_n_23_14),.A2(frontend_0_n_23_15),.ZN(frontend_0_n_23_16));
	OAI22_X1_LVT frontend_0i_23_17 (.A1(frontend_0_n_23_8),.A2(frontend_0_n_23_16),.B1(frontend_0_n_23_15),.B2(frontend_0_n_23_13),.ZN(frontend_0_n_18));
	NOR4_X1_LVT frontend_0i_41_0 (.A1(fe_mdb_in[0]),.A2(fe_mdb_in[1]),.A3(fe_mdb_in[2]),.A4(fe_mdb_in[3]),.ZN(frontend_0_n_48));
	AOI21_X1_LVT frontend_0i_44_0 (.A(frontend_0_n_49),.B1(frontend_0_n_18),.B2(frontend_0_n_48),.ZN(frontend_0_n_44_0));
	INV_X1_LVT frontend_0i_6_0 (.A(frontend_0_i_state[1]),.ZN(frontend_0_n_6_0));
	NOR3_X1_LVT frontend_0i_6_1 (.A1(frontend_0_n_6_0),.A2(frontend_0_i_state[0]),.A3(frontend_0_i_state[2]),.ZN(frontend_0_n_4));
	OR2_X1_LVT frontend_0i_61_0 (.A1(frontend_0_n_67),.A2(exec_done),.ZN(frontend_0_n_73));
	AND2_X1_LVT frontend_0i_62_0 (.A1(frontend_0_n_4),.A2(frontend_0_n_73),.ZN(decode_noirq));
	OR2_X1_LVT frontend_0i_63_0 (.A1(decode_noirq),.A2(frontend_0_irq_detect),.ZN(frontend_0_decode));
	INV_X1_LVT frontend_0i_44_1 (.A(frontend_0_decode),.ZN(frontend_0_n_44_1));
	NOR2_X1_LVT frontend_0i_44_2 (.A1(frontend_0_n_44_0),.A2(frontend_0_n_44_1),.ZN(frontend_0_n_51));
	INV_X1_LVT frontend_0i_45_0 (.A(frontend_0_n_51),.ZN(frontend_0_n_45_0));
	NAND3_X1_LVT frontend_0i_45_1 (.A1(frontend_0_n_45_0),.A2(e_state[2]),.A3(e_state[3]),.ZN(frontend_0_n_45_1));
	NOR3_X1_LVT frontend_0i_45_2 (.A1(frontend_0_n_45_1),.A2(e_state[0]),.A3(e_state[1]),.ZN(frontend_0_n_45_2));
	OR2_X1_LVT frontend_0i_45_3 (.A1(frontend_0_n_45_2),.A2(frontend_0_n_51),.ZN(frontend_0_n_52));
	CLKGATETST_X1_LVT frontend_0clk_gate_exec_jmp_reg (.CK(cpu_mclk),.E(frontend_0_n_52),.SE(1'b0),.GCK(frontend_0_n_50));
	DFFR_X1_LVT frontend_0exec_jmp_reg (.D(frontend_0_n_51),.RN(frontend_0_n_91),.CK(frontend_0_n_50),.Q(frontend_0_exec_jmp),.QN());
	NOR2_X1_LVT frontend_0i_59_0 (.A1(frontend_0_exec_dst_wr),.A2(frontend_0_exec_jmp),.ZN(frontend_0_n_59_0));
	AND2_X1_LVT frontend_0i_9_0 (.A1(frontend_0_n_10),.A2(frontend_0_n_9),.ZN(frontend_0_n_11));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_type_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_43));
	DFFR_X1_LVT frontend_0inst_type_reg___05F05b0___05F05d (.D(frontend_0_n_11),.RN(frontend_0_n_91),.CK(frontend_0_n_43),.Q(inst_type[0]),.QN());
	INV_X1_LVT frontend_0i_58_4 (.A(e_state[1]),.ZN(frontend_0_n_58_3));
	INV_X1_LVT frontend_0i_58_2 (.A(e_state[2]),.ZN(frontend_0_n_58_2));
	NOR4_X1_LVT frontend_0i_58_5 (.A1(frontend_0_n_58_3),.A2(frontend_0_n_58_2),.A3(e_state[0]),.A4(e_state[3]),.ZN(frontend_0_n_68));
	AND2_X1_LVT frontend_0i_37_0 (.A1(inst_type[0]),.A2(frontend_0_n_68),.ZN(frontend_0_n_45));
	INV_X1_LVT frontend_0i_58_1 (.A(e_state[0]),.ZN(frontend_0_n_58_1));
	NOR4_X1_LVT frontend_0i_58_6 (.A1(frontend_0_n_58_2),.A2(frontend_0_n_58_1),.A3(frontend_0_n_58_3),.A4(e_state[3]),.ZN(frontend_0_n_69));
	NOR4_X1_LVT frontend_0i_58_7 (.A1(frontend_0_n_58_3),.A2(frontend_0_n_58_0),.A3(e_state[0]),.A4(e_state[2]),.ZN(frontend_0_n_70));
	OR2_X1_LVT frontend_0i_38_0 (.A1(frontend_0_n_69),.A2(frontend_0_n_70),.ZN(frontend_0_n_46));
	INV_X1_LVT frontend_0i_39_1 (.A(frontend_0_n_46),.ZN(frontend_0_n_39_1));
	INV_X1_LVT frontend_0i_39_0 (.A(frontend_0_n_45),.ZN(frontend_0_n_39_0));
	NAND2_X1_LVT frontend_0i_39_2 (.A1(frontend_0_n_39_1),.A2(frontend_0_n_39_0),.ZN(frontend_0_n_47));
	CLKGATETST_X1_LVT frontend_0clk_gate_exec_src_wr_reg (.CK(cpu_mclk),.E(frontend_0_n_47),.SE(1'b0),.GCK(frontend_0_n_44));
	DFFR_X1_LVT frontend_0exec_src_wr_reg (.D(frontend_0_n_45),.RN(frontend_0_n_91),.CK(frontend_0_n_44),.Q(frontend_0_exec_src_wr),.QN());
	NAND3_X1_LVT frontend_0i_59_1 (.A1(frontend_0_n_59_0),.A2(frontend_0_exec_src_wr),.A3(frontend_0_n_69),.ZN(frontend_0_n_59_1));
	INV_X1_LVT frontend_0i_59_2 (.A(frontend_0_exec_src_wr),.ZN(frontend_0_n_59_2));
	NOR4_X1_LVT frontend_0i_58_9 (.A1(frontend_0_n_58_0),.A2(frontend_0_n_58_1),.A3(frontend_0_n_58_3),.A4(e_state[2]),.ZN(frontend_0_n_72));
	NAND3_X1_LVT frontend_0i_59_3 (.A1(frontend_0_n_59_0),.A2(frontend_0_n_59_2),.A3(frontend_0_n_72),.ZN(frontend_0_n_59_3));
	INV_X1_LVT frontend_0i_59_4 (.A(frontend_0_exec_jmp),.ZN(frontend_0_n_59_4));
	NAND3_X1_LVT frontend_0i_59_5 (.A1(frontend_0_n_59_4),.A2(frontend_0_exec_dst_wr),.A3(frontend_0_n_70),.ZN(frontend_0_n_59_5));
	NOR4_X1_LVT frontend_0i_58_8 (.A1(frontend_0_n_58_2),.A2(frontend_0_n_58_0),.A3(e_state[0]),.A4(e_state[1]),.ZN(frontend_0_n_71));
	NAND2_X1_LVT frontend_0i_59_6 (.A1(frontend_0_n_71),.A2(frontend_0_exec_jmp),.ZN(frontend_0_n_59_6));
	NAND4_X1_LVT frontend_0i_59_7 (.A1(frontend_0_n_59_1),.A2(frontend_0_n_59_3),.A3(frontend_0_n_59_5),.A4(frontend_0_n_59_6),.ZN(exec_done));
	OAI21_X1_LVT frontend_0i_60_0 (.A(frontend_0_n_3),.B1(frontend_0_n_5),.B2(exec_done),.ZN(frontend_0_n_60_0));
	INV_X1_LVT frontend_0i_60_1 (.A(frontend_0_n_60_0),.ZN(frontend_0_irq_detect));
	INV_X1_LVT frontend_0i_27_0 (.A(frontend_0_irq_detect),.ZN(frontend_0_n_27_0));
	NAND2_X1_LVT frontend_0i_27_9 (.A1(frontend_0_n_27_1),.A2(frontend_0_n_27_0),.ZN(frontend_0_inst_so_nxt[7]));
	AND2_X1_LVT frontend_0i_49_3 (.A1(frontend_0_n_1),.A2(frontend_0_inst_so_nxt[7]),.ZN(frontend_0_n_56));
	NOR2_X1_LVT frontend_0i_50_0 (.A1(frontend_0_n_55),.A2(frontend_0_n_56),.ZN(frontend_0_n_50_0));
	INV_X1_LVT frontend_0i_50_1 (.A(frontend_0_n_50_0),.ZN(frontend_0_n_50_1));
	NOR2_X1_LVT frontend_0i_50_2 (.A1(frontend_0_n_50_1),.A2(cpuoff),.ZN(frontend_0_n_50_2));
	INV_X1_LVT frontend_0i_50_3 (.A(frontend_0_n_50_2),.ZN(frontend_0_n_50_3));
	INV_X1_LVT frontend_0i_10_0 (.A(frontend_0_n_11),.ZN(frontend_0_n_10_0));
	AOI22_X1_LVT frontend_0i_10_1 (.A1(frontend_0_n_10_0),.A2(fe_mdb_in[8]),.B1(fe_mdb_in[0]),.B2(frontend_0_n_11),.ZN(frontend_0_n_10_1));
	INV_X1_LVT frontend_0i_10_2 (.A(frontend_0_n_10_1),.ZN(frontend_0_src_reg[0]));
	AOI22_X1_LVT frontend_0i_10_3 (.A1(frontend_0_n_10_0),.A2(fe_mdb_in[9]),.B1(frontend_0_n_11),.B2(fe_mdb_in[1]),.ZN(frontend_0_n_10_2));
	INV_X1_LVT frontend_0i_10_4 (.A(frontend_0_n_10_2),.ZN(frontend_0_src_reg[1]));
	AOI22_X1_LVT frontend_0i_10_5 (.A1(frontend_0_n_10_0),.A2(fe_mdb_in[10]),.B1(frontend_0_n_11),.B2(fe_mdb_in[2]),.ZN(frontend_0_n_10_3));
	INV_X1_LVT frontend_0i_10_6 (.A(frontend_0_n_10_3),.ZN(frontend_0_src_reg[2]));
	AOI22_X1_LVT frontend_0i_10_7 (.A1(frontend_0_n_10_0),.A2(fe_mdb_in[11]),.B1(frontend_0_n_11),.B2(fe_mdb_in[3]),.ZN(frontend_0_n_10_4));
	INV_X1_LVT frontend_0i_10_8 (.A(frontend_0_n_10_4),.ZN(frontend_0_src_reg[3]));
	NOR4_X1_LVT frontend_0i_12_12 (.A1(frontend_0_src_reg[0]),.A2(frontend_0_src_reg[1]),.A3(frontend_0_src_reg[2]),.A4(frontend_0_src_reg[3]),.ZN(frontend_0_n_12_11));
	INV_X1_LVT frontend_0i_12_16 (.A(frontend_0_n_12_11),.ZN(frontend_0_n_12_12));
	INV_X1_LVT frontend_0i_12_6 (.A(frontend_0_src_reg[0]),.ZN(frontend_0_n_12_6));
	INV_X1_LVT frontend_0i_12_7 (.A(frontend_0_src_reg[1]),.ZN(frontend_0_n_12_7));
	NOR4_X1_LVT frontend_0i_12_8 (.A1(frontend_0_n_12_6),.A2(frontend_0_n_12_7),.A3(frontend_0_src_reg[2]),.A4(frontend_0_src_reg[3]),.ZN(frontend_0_n_12_8));
	OR2_X1_LVT frontend_0i_12_9 (.A1(frontend_0_n_12_8),.A2(frontend_0_inst_type_nxt),.ZN(frontend_0_n_12_9));
	NOR4_X1_LVT frontend_0i_12_11 (.A1(frontend_0_n_12_7),.A2(frontend_0_src_reg[0]),.A3(frontend_0_src_reg[2]),.A4(frontend_0_src_reg[3]),.ZN(frontend_0_n_12_10));
	INV_X1_LVT frontend_0i_12_1 (.A(fe_mdb_in[5]),.ZN(frontend_0_n_12_1));
	NAND2_X1_LVT frontend_0i_12_3 (.A1(frontend_0_n_12_1),.A2(fe_mdb_in[4]),.ZN(frontend_0_n_12_3));
	NOR4_X1_LVT frontend_0i_12_17 (.A1(frontend_0_n_12_12),.A2(frontend_0_n_12_9),.A3(frontend_0_n_12_10),.A4(frontend_0_n_12_3),.ZN(frontend_0_inst_as_nxt[4]));
	INV_X1_LVT frontend_0i_12_19 (.A(frontend_0_n_12_10),.ZN(frontend_0_n_12_13));
	NOR3_X1_LVT frontend_0i_12_20 (.A1(frontend_0_n_12_13),.A2(frontend_0_n_12_9),.A3(frontend_0_n_12_3),.ZN(frontend_0_inst_as_nxt[6]));
	NOR4_X1_LVT frontend_0i_12_13 (.A1(frontend_0_n_12_9),.A2(frontend_0_n_12_10),.A3(frontend_0_n_12_3),.A4(frontend_0_n_12_11),.ZN(frontend_0_inst_as_nxt[1]));
	OR3_X1_LVT frontend_0i_48_0 (.A1(frontend_0_inst_as_nxt[4]),.A2(frontend_0_inst_as_nxt[6]),.A3(frontend_0_inst_as_nxt[1]),.ZN(frontend_0_src_acalc_pre));
	NOR2_X1_LVT frontend_0i_50_4 (.A1(frontend_0_n_50_3),.A2(frontend_0_src_acalc_pre),.ZN(frontend_0_n_50_4));
	OR2_X1_LVT frontend_0i_12_2 (.A1(frontend_0_n_12_1),.A2(fe_mdb_in[4]),.ZN(frontend_0_n_12_2));
	NOR3_X1_LVT frontend_0i_12_14 (.A1(frontend_0_n_12_9),.A2(frontend_0_n_12_10),.A3(frontend_0_n_12_2),.ZN(frontend_0_inst_as_nxt[2]));
	NAND2_X1_LVT frontend_0i_12_4 (.A1(fe_mdb_in[4]),.A2(fe_mdb_in[5]),.ZN(frontend_0_n_12_4));
	NOR4_X1_LVT frontend_0i_12_15 (.A1(frontend_0_n_12_9),.A2(frontend_0_n_12_10),.A3(frontend_0_n_12_11),.A4(frontend_0_n_12_4),.ZN(frontend_0_inst_as_nxt[3]));
	NOR4_X1_LVT frontend_0i_12_18 (.A1(frontend_0_n_12_12),.A2(frontend_0_n_12_9),.A3(frontend_0_n_12_10),.A4(frontend_0_n_12_4),.ZN(frontend_0_inst_as_nxt[5]));
	OR4_X1_LVT frontend_0i_49_1 (.A1(frontend_0_inst_as_nxt[2]),.A2(frontend_0_inst_as_nxt[3]),.A3(frontend_0_inst_as_nxt[5]),.A4(frontend_0_inst_so_nxt[6]),.ZN(frontend_0_n_54));
	INV_X1_LVT frontend_0i_50_5 (.A(frontend_0_n_54),.ZN(frontend_0_n_50_5));
	NAND2_X1_LVT frontend_0i_50_6 (.A1(frontend_0_n_50_4),.A2(frontend_0_n_50_5),.ZN(frontend_0_n_50_6));
	NOR2_X1_LVT frontend_0i_23_19 (.A1(frontend_0_n_23_3),.A2(frontend_0_n_23_16),.ZN(frontend_0_n_20));
	NOR3_X1_LVT frontend_0i_23_18 (.A1(frontend_0_n_23_16),.A2(frontend_0_n_23_6),.A3(frontend_0_n_23_0),.ZN(frontend_0_n_19));
	INV_X1_LVT frontend_0i_23_20 (.A(frontend_0_n_17),.ZN(frontend_0_n_23_17));
	NOR2_X1_LVT frontend_0i_23_21 (.A1(frontend_0_n_23_12),.A2(frontend_0_n_23_17),.ZN(frontend_0_inst_ad_nxt));
	OR3_X1_LVT frontend_0i_47_0 (.A1(frontend_0_n_20),.A2(frontend_0_n_19),.A3(frontend_0_inst_ad_nxt),.ZN(frontend_0_dst_acalc_pre));
	NOR2_X1_LVT frontend_0i_50_7 (.A1(frontend_0_n_50_6),.A2(frontend_0_dst_acalc_pre),.ZN(frontend_0_n_50_7));
	INV_X1_LVT frontend_0i_25_1 (.A(fe_mdb_in[8]),.ZN(frontend_0_n_25_1));
	NAND2_X1_LVT frontend_0i_25_2 (.A1(frontend_0_n_25_0),.A2(frontend_0_n_25_1),.ZN(frontend_0_n_25_2));
	NOR2_X1_LVT frontend_0i_25_11 (.A1(frontend_0_n_25_2),.A2(frontend_0_n_25_6),.ZN(frontend_0_n_26));
	AND2_X1_LVT frontend_0i_26_4 (.A1(frontend_0_n_10),.A2(frontend_0_n_26),.ZN(frontend_0_n_34));
	AND2_X1_LVT frontend_0i_27_5 (.A1(frontend_0_n_27_0),.A2(frontend_0_n_34),.ZN(frontend_0_inst_so_nxt[4]));
	NAND2_X1_LVT frontend_0i_25_3 (.A1(fe_mdb_in[7]),.A2(frontend_0_n_25_1),.ZN(frontend_0_n_25_3));
	NOR2_X1_LVT frontend_0i_25_12 (.A1(frontend_0_n_25_3),.A2(frontend_0_n_25_6),.ZN(frontend_0_n_27));
	AND2_X1_LVT frontend_0i_26_5 (.A1(frontend_0_n_10),.A2(frontend_0_n_27),.ZN(frontend_0_n_35));
	AND2_X1_LVT frontend_0i_27_6 (.A1(frontend_0_n_27_0),.A2(frontend_0_n_35),.ZN(frontend_0_inst_so_nxt[5]));
	OR2_X1_LVT frontend_0i_49_0 (.A1(frontend_0_inst_so_nxt[4]),.A2(frontend_0_inst_so_nxt[5]),.ZN(frontend_0_n_53));
	INV_X1_LVT frontend_0i_50_8 (.A(frontend_0_n_53),.ZN(frontend_0_n_50_8));
	NAND2_X1_LVT frontend_0i_50_9 (.A1(frontend_0_n_50_7),.A2(frontend_0_n_50_8),.ZN(frontend_0_n_50_9));
	NAND2_X1_LVT frontend_0i_50_17 (.A1(frontend_0_n_50_4),.A2(frontend_0_n_54),.ZN(frontend_0_n_50_16));
	INV_X1_LVT frontend_0i_50_12 (.A(frontend_0_n_56),.ZN(frontend_0_n_50_12));
	NAND3_X1_LVT frontend_0i_50_18 (.A1(frontend_0_n_50_9),.A2(frontend_0_n_50_16),.A3(frontend_0_n_50_12),.ZN(frontend_0_n_58));
	AND2_X1_LVT frontend_0i_55_36 (.A1(frontend_0_n_55_6),.A2(frontend_0_n_58),.ZN(frontend_0_n_55_35));
	NOR4_X1_LVT frontend_0i_55_18 (.A1(e_state[0]),.A2(e_state[1]),.A3(e_state[2]),.A4(e_state[3]),.ZN(frontend_0_n_55_18));
	NAND4_X1_LVT frontend_0i_55_23 (.A1(frontend_0_n_55_1),.A2(frontend_0_n_55_10),.A3(e_state[0]),.A4(e_state[3]),.ZN(frontend_0_n_55_23));
	INV_X1_LVT frontend_0i_55_37 (.A(frontend_0_n_55_23),.ZN(frontend_0_n_55_36));
	NOR4_X1_LVT frontend_0i_55_38 (.A1(frontend_0_n_55_35),.A2(frontend_0_n_55_18),.A3(frontend_0_n_55_21),.A4(frontend_0_n_55_36),.ZN(frontend_0_n_55_37));
	NOR4_X1_LVT frontend_0i_55_30 (.A1(frontend_0_n_55_0),.A2(frontend_0_n_55_10),.A3(e_state[1]),.A4(e_state[3]),.ZN(frontend_0_n_55_30));
	NOR3_X1_LVT frontend_0i_6_5 (.A1(frontend_0_n_6_0),.A2(frontend_0_n_6_2),.A3(frontend_0_i_state[2]),.ZN(frontend_0_n_6));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_as_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_12));
	DFFR_X1_LVT frontend_0inst_as_reg___05F05b6___05F05d (.D(frontend_0_inst_as_nxt[6]),.RN(frontend_0_n_91),.CK(frontend_0_n_12),.Q(inst_as[6]),.QN());
	DFFR_X1_LVT frontend_0inst_as_reg___05F05b1___05F05d (.D(frontend_0_inst_as_nxt[1]),.RN(frontend_0_n_91),.CK(frontend_0_n_12),.Q(inst_as[1]),.QN());
	DFFR_X1_LVT frontend_0inst_as_reg___05F05b5___05F05d (.D(frontend_0_inst_as_nxt[5]),.RN(frontend_0_n_91),.CK(frontend_0_n_12),.Q(inst_as[5]),.QN());
	DFFR_X1_LVT frontend_0inst_as_reg___05F05b4___05F05d (.D(frontend_0_inst_as_nxt[4]),.RN(frontend_0_n_91),.CK(frontend_0_n_12),.Q(inst_as[4]),.QN());
	OR4_X1_LVT frontend_0i_15_0 (.A1(inst_as[6]),.A2(inst_as[1]),.A3(inst_as[5]),.A4(inst_as[4]),.ZN(frontend_0_is_sext));
	AND2_X1_LVT frontend_0i_30_0 (.A1(frontend_0_n_6),.A2(frontend_0_is_sext),.ZN(frontend_0_inst_sext_rdy));
	NAND2_X1_LVT frontend_0i_55_39 (.A1(frontend_0_n_55_30),.A2(frontend_0_inst_sext_rdy),.ZN(frontend_0_n_55_38));
	INV_X1_LVT frontend_0i_55_4 (.A(e_state[3]),.ZN(frontend_0_n_55_4));
	NAND4_X1_LVT frontend_0i_55_32 (.A1(frontend_0_n_55_0),.A2(frontend_0_n_55_4),.A3(e_state[1]),.A4(e_state[2]),.ZN(frontend_0_n_55_32));
	INV_X1_LVT frontend_0i_55_33 (.A(frontend_0_n_55_32),.ZN(frontend_0_n_55_33));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_so_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_38));
	DFFR_X1_LVT frontend_0inst_so_reg___05F05b6___05F05d (.D(frontend_0_inst_so_nxt[6]),.RN(frontend_0_n_91),.CK(frontend_0_n_38),.Q(inst_so[6]),.QN());
	DFFR_X1_LVT frontend_0inst_so_reg___05F05b4___05F05d (.D(frontend_0_inst_so_nxt[4]),.RN(frontend_0_n_91),.CK(frontend_0_n_38),.Q(inst_so[4]),.QN());
	DFFR_X1_LVT frontend_0inst_so_reg___05F05b5___05F05d (.D(frontend_0_inst_so_nxt[5]),.RN(frontend_0_n_91),.CK(frontend_0_n_38),.Q(inst_so[5]),.QN());
	OR2_X1_LVT frontend_0i_29_0 (.A1(inst_so[4]),.A2(inst_so[5]),.ZN(frontend_0_n_39));
	OR2_X1_LVT frontend_0i_52_0 (.A1(inst_so[6]),.A2(frontend_0_n_39),.ZN(frontend_0_n_62));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_ad_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_21));
	DFFR_X1_LVT frontend_0inst_ad_reg___05F05b4___05F05d (.D(frontend_0_n_20),.RN(frontend_0_n_91),.CK(frontend_0_n_21),.Q(inst_ad[4]),.QN());
	DFFR_X1_LVT frontend_0inst_ad_reg___05F05b1___05F05d (.D(frontend_0_n_19),.RN(frontend_0_n_91),.CK(frontend_0_n_21),.Q(inst_ad[1]),.QN());
	DFFR_X1_LVT frontend_0inst_ad_reg___05F05b6___05F05d (.D(frontend_0_inst_ad_nxt),.RN(frontend_0_n_91),.CK(frontend_0_n_21),.Q(inst_ad[6]),.QN());
	OR3_X1_LVT frontend_0i_52_1 (.A1(inst_ad[4]),.A2(inst_ad[1]),.A3(inst_ad[6]),.ZN(frontend_0_n_63));
	NOR2_X1_LVT frontend_0i_53_0 (.A1(frontend_0_n_62),.A2(frontend_0_n_63),.ZN(frontend_0_n_64));
	NAND2_X1_LVT frontend_0i_55_40 (.A1(frontend_0_n_55_33),.A2(frontend_0_n_64),.ZN(frontend_0_n_55_39));
	NAND4_X1_LVT frontend_0i_55_11 (.A1(frontend_0_n_55_10),.A2(e_state[0]),.A3(e_state[1]),.A4(e_state[3]),.ZN(frontend_0_n_55_11));
	INV_X1_LVT frontend_0i_55_41 (.A(frontend_0_n_55_11),.ZN(frontend_0_n_55_40));
	NOR2_X1_LVT frontend_0i_55_12 (.A1(frontend_0_exec_jmp),.A2(frontend_0_exec_dst_wr),.ZN(frontend_0_n_55_12));
	NAND2_X1_LVT frontend_0i_55_16 (.A1(frontend_0_n_55_12),.A2(frontend_0_exec_src_wr),.ZN(frontend_0_n_55_16));
	INV_X1_LVT frontend_0i_55_13 (.A(frontend_0_n_55_12),.ZN(frontend_0_n_55_13));
	NOR2_X1_LVT frontend_0i_55_14 (.A1(frontend_0_n_55_13),.A2(frontend_0_exec_src_wr),.ZN(frontend_0_n_55_14));
	INV_X1_LVT frontend_0i_55_43 (.A(frontend_0_n_55_14),.ZN(frontend_0_n_55_42));
	INV_X1_LVT frontend_0i_55_44 (.A(frontend_0_n_58),.ZN(frontend_0_n_55_43));
	OAI211_X1_LVT frontend_0i_55_45 (.A(frontend_0_n_55_16),.B(frontend_0_n_55_41),.C1(frontend_0_n_55_42),.C2(frontend_0_n_55_43),.ZN(frontend_0_n_55_44));
	NAND2_X1_LVT frontend_0i_55_46 (.A1(frontend_0_n_55_40),.A2(frontend_0_n_55_44),.ZN(frontend_0_n_55_45));
	AND4_X1_LVT frontend_0i_55_47 (.A1(frontend_0_n_55_37),.A2(frontend_0_n_55_38),.A3(frontend_0_n_55_39),.A4(frontend_0_n_55_45),.ZN(frontend_0_n_55_46));
	NAND4_X1_LVT frontend_0i_55_26 (.A1(frontend_0_n_55_0),.A2(frontend_0_n_55_10),.A3(e_state[1]),.A4(e_state[3]),.ZN(frontend_0_n_55_26));
	INV_X1_LVT frontend_0i_55_27 (.A(frontend_0_n_55_26),.ZN(frontend_0_n_55_27));
	INV_X1_LVT frontend_0i_55_28 (.A(frontend_0_exec_jmp),.ZN(frontend_0_n_55_28));
	NAND3_X1_LVT frontend_0i_55_48 (.A1(frontend_0_n_55_27),.A2(frontend_0_n_55_28),.A3(frontend_0_n_58),.ZN(frontend_0_n_55_47));
	NAND4_X1_LVT frontend_0i_55_3 (.A1(frontend_0_n_55_1),.A2(e_state[0]),.A3(e_state[2]),.A4(e_state[3]),.ZN(frontend_0_n_55_3));
	NAND4_X1_LVT frontend_0i_55_5 (.A1(frontend_0_n_55_4),.A2(e_state[0]),.A3(e_state[1]),.A4(e_state[2]),.ZN(frontend_0_n_55_5));
	AND4_X1_LVT frontend_0i_55_49 (.A1(frontend_0_n_55_26),.A2(frontend_0_n_55_3),.A3(frontend_0_n_55_11),.A4(frontend_0_n_55_5),.ZN(frontend_0_n_55_48));
	NAND4_X1_LVT frontend_0i_55_50 (.A1(frontend_0_n_55_48),.A2(frontend_0_n_55_32),.A3(frontend_0_n_55_23),.A4(frontend_0_n_55_2),.ZN(frontend_0_n_55_49));
	NOR4_X1_LVT frontend_0i_55_8 (.A1(frontend_0_n_55_4),.A2(e_state[0]),.A3(e_state[1]),.A4(e_state[2]),.ZN(frontend_0_n_55_8));
	NOR4_X1_LVT frontend_0i_55_51 (.A1(frontend_0_n_55_0),.A2(frontend_0_n_55_1),.A3(e_state[2]),.A4(e_state[3]),.ZN(frontend_0_n_55_50));
	NOR4_X1_LVT frontend_0i_55_52 (.A1(frontend_0_n_55_49),.A2(frontend_0_n_55_8),.A3(frontend_0_n_55_50),.A4(frontend_0_n_55_30),.ZN(frontend_0_n_55_51));
	NAND4_X1_LVT frontend_0i_55_20 (.A1(frontend_0_n_55_0),.A2(frontend_0_n_55_10),.A3(frontend_0_n_55_4),.A4(e_state[1]),.ZN(frontend_0_n_55_20));
	NAND4_X1_LVT frontend_0i_55_53 (.A1(frontend_0_n_55_1),.A2(frontend_0_n_55_10),.A3(frontend_0_n_55_4),.A4(e_state[0]),.ZN(frontend_0_n_55_52));
	INV_X1_LVT frontend_0i_55_22 (.A(frontend_0_n_55_21),.ZN(frontend_0_n_55_22));
	NAND4_X1_LVT frontend_0i_55_54 (.A1(frontend_0_n_55_51),.A2(frontend_0_n_55_20),.A3(frontend_0_n_55_52),.A4(frontend_0_n_55_22),.ZN(frontend_0_n_55_53));
	OAI211_X1_LVT frontend_0i_55_55 (.A(frontend_0_n_55_46),.B(frontend_0_n_55_47),.C1(frontend_0_n_55_53),.C2(frontend_0_n_55_18),.ZN(frontend_0_e_state_nxt_reg[1]));
	DFFR_X1_LVT frontend_0e_state_reg___05F05b1___05F05d (.D(frontend_0_e_state_nxt_reg[1]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(e_state[1]),.QN());
	INV_X1_LVT frontend_0i_55_1 (.A(e_state[1]),.ZN(frontend_0_n_55_1));
	NAND4_X1_LVT frontend_0i_55_2 (.A1(frontend_0_n_55_0),.A2(frontend_0_n_55_1),.A3(e_state[2]),.A4(e_state[3]),.ZN(frontend_0_n_55_2));
	NAND3_X1_LVT frontend_0i_55_6 (.A1(frontend_0_n_55_2),.A2(frontend_0_n_55_3),.A3(frontend_0_n_55_5),.ZN(frontend_0_n_55_6));
	NAND2_X1_LVT frontend_0i_50_10 (.A1(frontend_0_n_50_2),.A2(frontend_0_src_acalc_pre),.ZN(frontend_0_n_50_10));
	NAND2_X1_LVT frontend_0i_50_11 (.A1(frontend_0_n_50_0),.A2(cpuoff),.ZN(frontend_0_n_50_11));
	NAND2_X1_LVT frontend_0i_50_13 (.A1(frontend_0_n_50_12),.A2(frontend_0_n_55),.ZN(frontend_0_n_50_13));
	AND4_X1_LVT frontend_0i_50_14 (.A1(frontend_0_n_50_9),.A2(frontend_0_n_50_10),.A3(frontend_0_n_50_11),.A4(frontend_0_n_50_13),.ZN(frontend_0_n_50_14));
	NAND2_X1_LVT frontend_0i_50_15 (.A1(frontend_0_n_50_7),.A2(frontend_0_n_53),.ZN(frontend_0_n_50_15));
	NAND2_X1_LVT frontend_0i_50_16 (.A1(frontend_0_n_50_14),.A2(frontend_0_n_50_15),.ZN(frontend_0_n_57));
	AND2_X1_LVT frontend_0i_55_7 (.A1(frontend_0_n_55_6),.A2(frontend_0_n_57),.ZN(frontend_0_n_55_7));
	INV_X1_LVT frontend_0i_16_0 (.A(frontend_0_n_6),.ZN(frontend_0_n_16_0));
	NOR2_X1_LVT frontend_0i_16_1 (.A1(frontend_0_n_16_0),.A2(frontend_0_is_sext),.ZN(frontend_0_n_13));
	NOR3_X1_LVT frontend_0i_6_6 (.A1(frontend_0_n_6_1),.A2(frontend_0_i_state[0]),.A3(frontend_0_i_state[1]),.ZN(frontend_0_n_7));
	OR2_X1_LVT frontend_0i_17_0 (.A1(frontend_0_n_13),.A2(frontend_0_n_7),.ZN(frontend_0_inst_dext_rdy));
	NAND2_X1_LVT frontend_0i_19_0 (.A1(e_state[0]),.A2(e_state[3]),.ZN(frontend_0_n_19_0));
	OR3_X1_LVT frontend_0i_19_1 (.A1(frontend_0_n_19_0),.A2(e_state[1]),.A3(e_state[2]),.ZN(frontend_0_n_19_1));
	AND2_X1_LVT frontend_0i_19_2 (.A1(frontend_0_n_19_1),.A2(frontend_0_inst_dext_rdy),.ZN(frontend_0_n_15));
	INV_X1_LVT frontend_0i_20_3 (.A(frontend_0_inst_dext_rdy),.ZN(frontend_0_n_20_3));
	NAND2_X1_LVT frontend_0i_20_0 (.A1(e_state[0]),.A2(e_state[3]),.ZN(frontend_0_n_20_0));
	NOR3_X1_LVT frontend_0i_20_1 (.A1(frontend_0_n_20_0),.A2(e_state[1]),.A3(e_state[2]),.ZN(frontend_0_n_20_1));
	INV_X1_LVT frontend_0i_20_2 (.A(frontend_0_n_20_1),.ZN(frontend_0_n_20_2));
	NAND2_X1_LVT frontend_0i_20_4 (.A1(frontend_0_n_20_3),.A2(frontend_0_n_20_2),.ZN(frontend_0_n_16));
	CLKGATETST_X1_LVT frontend_0clk_gate_exec_dext_rdy_reg (.CK(cpu_mclk),.E(frontend_0_n_16),.SE(1'b0),.GCK(frontend_0_n_14));
	DFFR_X1_LVT frontend_0exec_dext_rdy_reg (.D(frontend_0_n_15),.RN(frontend_0_n_91),.CK(frontend_0_n_14),.Q(frontend_0_exec_dext_rdy),.QN());
	OR2_X1_LVT frontend_0i_51_0 (.A1(frontend_0_inst_dext_rdy),.A2(frontend_0_exec_dext_rdy),.ZN(frontend_0_n_61));
	AND2_X1_LVT frontend_0i_55_9 (.A1(frontend_0_n_55_8),.A2(frontend_0_n_61),.ZN(frontend_0_n_55_9));
	NAND2_X1_LVT frontend_0i_55_15 (.A1(frontend_0_n_55_14),.A2(frontend_0_n_57),.ZN(frontend_0_n_55_15));
	AOI21_X1_LVT frontend_0i_55_17 (.A(frontend_0_n_55_11),.B1(frontend_0_n_55_15),.B2(frontend_0_n_55_16),.ZN(frontend_0_n_55_17));
	INV_X1_LVT frontend_0i_55_19 (.A(frontend_0_n_55_18),.ZN(frontend_0_n_55_19));
	NAND4_X1_LVT frontend_0i_55_24 (.A1(frontend_0_n_55_19),.A2(frontend_0_n_55_20),.A3(frontend_0_n_55_22),.A4(frontend_0_n_55_23),.ZN(frontend_0_n_55_24));
	NOR4_X1_LVT frontend_0i_55_25 (.A1(frontend_0_n_55_7),.A2(frontend_0_n_55_9),.A3(frontend_0_n_55_17),.A4(frontend_0_n_55_24),.ZN(frontend_0_n_55_25));
	NAND3_X1_LVT frontend_0i_55_29 (.A1(frontend_0_n_55_27),.A2(frontend_0_n_55_28),.A3(frontend_0_n_57),.ZN(frontend_0_n_55_29));
	INV_X1_LVT frontend_0i_54_0 (.A(frontend_0_inst_sext_rdy),.ZN(frontend_0_n_66));
	NAND2_X1_LVT frontend_0i_55_31 (.A1(frontend_0_n_55_30),.A2(frontend_0_n_66),.ZN(frontend_0_n_55_31));
	INV_X1_LVT frontend_0i_53_1 (.A(frontend_0_n_64),.ZN(frontend_0_n_53_0));
	INV_X1_LVT frontend_0i_53_2 (.A(frontend_0_n_62),.ZN(frontend_0_n_53_1));
	OAI21_X1_LVT frontend_0i_53_3 (.A(frontend_0_n_53_0),.B1(frontend_0_n_53_1),.B2(frontend_0_n_63),.ZN(frontend_0_n_65));
	NAND2_X1_LVT frontend_0i_55_34 (.A1(frontend_0_n_55_33),.A2(frontend_0_n_65),.ZN(frontend_0_n_55_34));
	NAND4_X1_LVT frontend_0i_55_35 (.A1(frontend_0_n_55_25),.A2(frontend_0_n_55_29),.A3(frontend_0_n_55_31),.A4(frontend_0_n_55_34),.ZN(frontend_0_e_state_nxt_reg[0]));
	DFFS_X1_LVT frontend_0e_state_reg___05F05b0___05F05d (.D(frontend_0_e_state_nxt_reg[0]),.SN(frontend_0_n_91),.CK(cpu_mclk),.Q(e_state[0]),.QN());
	NAND2_X1_LVT frontend_0i_32_0 (.A1(e_state[0]),.A2(e_state[3]),.ZN(frontend_0_n_32_0));
	NOR3_X1_LVT frontend_0i_32_1 (.A1(frontend_0_n_32_0),.A2(e_state[1]),.A3(e_state[2]),.ZN(frontend_0_n_41));
	INV_X1_LVT frontend_0i_33_0 (.A(e_state[1]),.ZN(frontend_0_n_33_0));
	INV_X1_LVT frontend_0i_33_1 (.A(e_state[2]),.ZN(frontend_0_n_33_1));
	NAND4_X1_LVT frontend_0i_33_2 (.A1(frontend_0_n_33_0),.A2(frontend_0_n_33_1),.A3(e_state[0]),.A4(e_state[3]),.ZN(frontend_0_n_33_2));
	INV_X1_LVT frontend_0i_33_3 (.A(e_state[0]),.ZN(frontend_0_n_33_3));
	NAND4_X1_LVT frontend_0i_33_4 (.A1(frontend_0_n_33_3),.A2(frontend_0_n_33_1),.A3(e_state[1]),.A4(e_state[3]),.ZN(frontend_0_n_33_4));
	NAND2_X1_LVT frontend_0i_33_5 (.A1(frontend_0_n_33_2),.A2(frontend_0_n_33_4),.ZN(frontend_0_n_42));
	CLKGATETST_X1_LVT frontend_0clk_gate_exec_dst_wr_reg (.CK(cpu_mclk),.E(frontend_0_n_42),.SE(1'b0),.GCK(frontend_0_n_40));
	DFFR_X1_LVT frontend_0exec_dst_wr_reg (.D(frontend_0_n_41),.RN(frontend_0_n_91),.CK(frontend_0_n_40),.Q(frontend_0_exec_dst_wr),.QN());
	INV_X1_LVT frontend_0i_55_42 (.A(frontend_0_exec_dst_wr),.ZN(frontend_0_n_55_41));
	NAND2_X1_LVT frontend_0i_55_56 (.A1(frontend_0_n_55_41),.A2(frontend_0_exec_jmp),.ZN(frontend_0_n_55_54));
	INV_X1_LVT frontend_0i_55_57 (.A(frontend_0_n_55_54),.ZN(frontend_0_n_55_55));
	INV_X1_LVT frontend_0i_55_58 (.A(frontend_0_n_55_16),.ZN(frontend_0_n_55_56));
	NAND4_X1_LVT frontend_0i_50_19 (.A1(frontend_0_n_50_16),.A2(frontend_0_n_50_10),.A3(frontend_0_n_50_11),.A4(frontend_0_n_50_13),.ZN(frontend_0_n_59));
	AOI211_X1_LVT frontend_0i_55_59 (.A(frontend_0_n_55_55),.B(frontend_0_n_55_56),.C1(frontend_0_n_55_14),.C2(frontend_0_n_59),.ZN(frontend_0_n_55_57));
	NOR2_X1_LVT frontend_0i_55_60 (.A1(frontend_0_n_55_57),.A2(frontend_0_n_55_11),.ZN(frontend_0_n_55_58));
	AND2_X1_LVT frontend_0i_55_61 (.A1(frontend_0_n_55_6),.A2(frontend_0_n_59),.ZN(frontend_0_n_55_59));
	NOR4_X1_LVT frontend_0i_55_62 (.A1(frontend_0_n_55_58),.A2(frontend_0_n_55_59),.A3(frontend_0_n_55_50),.A4(frontend_0_n_55_30),.ZN(frontend_0_n_55_60));
	NOR2_X1_LVT frontend_0i_55_72 (.A1(frontend_0_n_59),.A2(frontend_0_exec_jmp),.ZN(frontend_0_n_55_68));
	OAI21_X1_LVT frontend_0i_55_63 (.A(frontend_0_n_55_60),.B1(frontend_0_n_55_26),.B2(frontend_0_n_55_68),.ZN(frontend_0_e_state_nxt_reg[2]));
	DFFR_X1_LVT frontend_0e_state_reg___05F05b2___05F05d (.D(frontend_0_e_state_nxt_reg[2]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(e_state[2]),.QN());
	INV_X1_LVT frontend_0i_55_10 (.A(e_state[2]),.ZN(frontend_0_n_55_10));
	NOR4_X1_LVT frontend_0i_55_21 (.A1(frontend_0_n_55_10),.A2(e_state[0]),.A3(e_state[1]),.A4(e_state[3]),.ZN(frontend_0_n_55_21));
	NOR4_X1_LVT frontend_0i_55_64 (.A1(frontend_0_n_55_21),.A2(frontend_0_n_55_36),.A3(frontend_0_n_55_33),.A4(frontend_0_n_55_8),.ZN(frontend_0_n_55_61));
	INV_X1_LVT frontend_0i_50_20 (.A(frontend_0_n_50_6),.ZN(frontend_0_n_50_17));
	NAND2_X1_LVT frontend_0i_50_21 (.A1(frontend_0_n_50_17),.A2(frontend_0_dst_acalc_pre),.ZN(frontend_0_n_50_18));
	AND4_X1_LVT frontend_0i_50_22 (.A1(frontend_0_n_50_9),.A2(frontend_0_n_50_18),.A3(frontend_0_n_50_11),.A4(frontend_0_n_50_13),.ZN(frontend_0_n_50_19));
	NAND2_X1_LVT frontend_0i_50_23 (.A1(frontend_0_n_50_19),.A2(frontend_0_n_50_15),.ZN(frontend_0_n_60));
	INV_X1_LVT frontend_0i_55_65 (.A(frontend_0_n_60),.ZN(frontend_0_n_55_62));
	NOR2_X1_LVT frontend_0i_55_66 (.A1(frontend_0_n_55_62),.A2(frontend_0_exec_jmp),.ZN(frontend_0_n_55_63));
	OAI21_X1_LVT frontend_0i_55_67 (.A(frontend_0_n_55_27),.B1(frontend_0_n_55_63),.B2(frontend_0_exec_jmp),.ZN(frontend_0_n_55_64));
	OAI211_X1_LVT frontend_0i_55_68 (.A(frontend_0_n_55_54),.B(frontend_0_n_55_41),.C1(frontend_0_n_55_42),.C2(frontend_0_n_55_62),.ZN(frontend_0_n_55_65));
	NAND2_X1_LVT frontend_0i_55_69 (.A1(frontend_0_n_55_40),.A2(frontend_0_n_55_65),.ZN(frontend_0_n_55_66));
	NAND2_X1_LVT frontend_0i_55_70 (.A1(frontend_0_n_55_6),.A2(frontend_0_n_60),.ZN(frontend_0_n_55_67));
	NAND4_X1_LVT frontend_0i_55_71 (.A1(frontend_0_n_55_61),.A2(frontend_0_n_55_64),.A3(frontend_0_n_55_66),.A4(frontend_0_n_55_67),.ZN(frontend_0_e_state_nxt_reg[3]));
	DFFR_X1_LVT frontend_0e_state_reg___05F05b3___05F05d (.D(frontend_0_e_state_nxt_reg[3]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(e_state[3]),.QN());
	INV_X1_LVT frontend_0i_58_0 (.A(e_state[3]),.ZN(frontend_0_n_58_0));
	NOR4_X1_LVT frontend_0i_58_3 (.A1(frontend_0_n_58_0),.A2(frontend_0_n_58_1),.A3(frontend_0_n_58_2),.A4(e_state[1]),.ZN(frontend_0_n_67));
	AND2_X1_LVT frontend_0i_72_0 (.A1(frontend_0_cpu_halt_req),.A2(frontend_0_n_67),.ZN(frontend_0_n_82));
	OAI21_X1_LVT frontend_0i_72_1 (.A(exec_done),.B1(frontend_0_cpu_halt_req),.B2(cpuoff),.ZN(frontend_0_n_72_0));
	INV_X1_LVT frontend_0i_72_2 (.A(frontend_0_n_72_0),.ZN(frontend_0_n_83));
	NOR2_X1_LVT frontend_0i_73_0 (.A1(frontend_0_n_82),.A2(frontend_0_n_83),.ZN(frontend_0_n_73_0));
	NOR2_X1_LVT frontend_0i_73_6 (.A1(frontend_0_n_73_0),.A2(frontend_0_irq_detect),.ZN(frontend_0_n_86));
	NOR3_X1_LVT frontend_0i_76_13 (.A1(frontend_0_n_76_5),.A2(frontend_0_n_76_2),.A3(frontend_0_i_state[2]),.ZN(frontend_0_n_76_12));
	INV_X1_LVT frontend_0i_71_0 (.A(pc_sw_wr),.ZN(frontend_0_n_71_0));
	INV_X1_LVT frontend_0i_64_0 (.A(frontend_0_dst_acalc_pre),.ZN(frontend_0_n_64_0));
	NOR2_X1_LVT frontend_0i_64_1 (.A1(frontend_0_n_64_0),.A2(frontend_0_n_11),.ZN(frontend_0_n_74));
	OR2_X1_LVT frontend_0i_65_0 (.A1(frontend_0_inst_as_nxt[5]),.A2(frontend_0_src_acalc_pre),.ZN(frontend_0_n_75));
	HA_X1_LVT frontend_0i_66_0 (.A(frontend_0_n_74),.B(frontend_0_n_75),.CO(frontend_0_inst_sz_nxt[1]),.S(frontend_0_inst_sz_nxt[0]));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_sz_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_76));
	DFFR_X1_LVT frontend_0inst_sz_reg___05F05b1___05F05d (.D(frontend_0_inst_sz_nxt[1]),.RN(frontend_0_n_91),.CK(frontend_0_n_76),.Q(frontend_0_inst_sz[1]),.QN());
	INV_X1_LVT frontend_0i_70_0 (.A(frontend_0_inst_sz[1]),.ZN(frontend_0_n_70_0));
	DFFR_X1_LVT frontend_0inst_sz_reg___05F05b0___05F05d (.D(frontend_0_inst_sz_nxt[0]),.RN(frontend_0_n_91),.CK(frontend_0_n_76),.Q(frontend_0_inst_sz[0]),.QN());
	NAND2_X1_LVT frontend_0i_70_1 (.A1(frontend_0_n_70_0),.A2(frontend_0_inst_sz[0]),.ZN(frontend_0_n_79));
	AND2_X1_LVT frontend_0i_71_1 (.A1(frontend_0_n_71_0),.A2(frontend_0_n_79),.ZN(frontend_0_n_80));
	AOI221_X1_LVT frontend_0i_76_16 (.A(frontend_0_n_76_4),.B1(frontend_0_n_76_6),.B2(frontend_0_n_86),.C1(frontend_0_n_76_12),.C2(frontend_0_n_80),.ZN(frontend_0_n_76_14));
	INV_X1_LVT frontend_0i_76_17 (.A(frontend_0_n_76_14),.ZN(frontend_0_i_state_nxt_reg[2]));
	DFFR_X1_LVT frontend_0i_state_reg___05F05b2___05F05d (.D(frontend_0_i_state_nxt_reg[2]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(frontend_0_i_state[2]),.QN());
	OAI33_X1_LVT frontend_0i_76_9 (.A1(frontend_0_n_76_2),.A2(frontend_0_i_state[1]),.A3(frontend_0_i_state[2]),.B1(frontend_0_n_76_1),.B2(frontend_0_i_state[0]),.B3(frontend_0_i_state[1]),.ZN(frontend_0_n_76_8));
	INV_X1_LVT frontend_0i_76_10 (.A(frontend_0_n_76_8),.ZN(frontend_0_n_76_9));
	INV_X1_LVT frontend_0i_75_1 (.A(frontend_0_n_87),.ZN(frontend_0_n_75_0));
	NOR2_X1_LVT frontend_0i_75_2 (.A1(frontend_0_n_75_0),.A2(frontend_0_n_88),.ZN(frontend_0_n_90));
	NAND2_X1_LVT frontend_0i_76_11 (.A1(frontend_0_n_76_3),.A2(frontend_0_n_90),.ZN(frontend_0_n_76_10));
	INV_X1_LVT frontend_0i_73_1 (.A(frontend_0_n_73_0),.ZN(frontend_0_n_73_1));
	NOR2_X1_LVT frontend_0i_73_5 (.A1(frontend_0_n_73_1),.A2(frontend_0_irq_detect),.ZN(frontend_0_n_85));
	NAND2_X1_LVT frontend_0i_76_12 (.A1(frontend_0_n_76_6),.A2(frontend_0_n_85),.ZN(frontend_0_n_76_11));
	INV_X1_LVT frontend_0i_71_2 (.A(frontend_0_n_80),.ZN(frontend_0_n_81));
	NAND2_X1_LVT frontend_0i_76_14 (.A1(frontend_0_n_76_12),.A2(frontend_0_n_81),.ZN(frontend_0_n_76_13));
	NAND4_X1_LVT frontend_0i_76_15 (.A1(frontend_0_n_76_9),.A2(frontend_0_n_76_10),.A3(frontend_0_n_76_11),.A4(frontend_0_n_76_13),.ZN(frontend_0_i_state_nxt_reg[1]));
	DFFR_X1_LVT frontend_0i_state_reg___05F05b1___05F05d (.D(frontend_0_i_state_nxt_reg[1]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(frontend_0_i_state[1]),.QN());
	NOR3_X1_LVT frontend_0i_76_0 (.A1(frontend_0_i_state[0]),.A2(frontend_0_i_state[1]),.A3(frontend_0_i_state[2]),.ZN(frontend_0_n_76_0));
	NOR2_X1_LVT frontend_0i_68_0 (.A1(exec_done),.A2(frontend_0_n_67),.ZN(frontend_0_n_77));
	OR2_X1_LVT frontend_0i_69_0 (.A1(frontend_0_inst_sz_nxt[0]),.A2(frontend_0_inst_sz_nxt[1]),.ZN(frontend_0_n_78));
	INV_X1_LVT frontend_0i_73_2 (.A(frontend_0_n_78),.ZN(frontend_0_n_73_2));
	OR4_X1_LVT frontend_0i_73_3 (.A1(frontend_0_n_73_1),.A2(frontend_0_n_77),.A3(pc_sw_wr),.A4(frontend_0_n_73_2),.ZN(frontend_0_n_73_3));
	AOI21_X1_LVT frontend_0i_73_4 (.A(frontend_0_irq_detect),.B1(frontend_0_n_73_3),.B2(frontend_0_n_73_0),.ZN(frontend_0_n_84));
	AOI211_X1_LVT frontend_0i_76_7 (.A(frontend_0_n_76_0),.B(frontend_0_n_76_4),.C1(frontend_0_n_76_6),.C2(frontend_0_n_84),.ZN(frontend_0_n_76_7));
	INV_X1_LVT frontend_0i_76_8 (.A(frontend_0_n_76_7),.ZN(frontend_0_i_state_nxt_reg[0]));
	NAND3_X1_LVT frontend_0i_80_0 (.A1(frontend_0_i_state_nxt_reg[0]),.A2(frontend_0_i_state_nxt_reg[2]),.A3(frontend_0_cpu_halt_req),.ZN(frontend_0_n_80_0));
	NOR2_X1_LVT frontend_0i_80_1 (.A1(frontend_0_n_80_0),.A2(frontend_0_i_state_nxt_reg[1]),.ZN(frontend_0_n_92));
	DFFR_X1_LVT frontend_0cpu_halt_st_reg (.D(frontend_0_n_92),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(cpu_halt_st),.QN());
	DFFR_X1_LVT frontend_0inst_ad_reg___05F05b7___05F05d (.D(1'b0),.RN(frontend_0_n_91),.CK(frontend_0_n_21),.Q(inst_ad[7]),.QN());
	DFFR_X1_LVT frontend_0inst_ad_reg___05F05b5___05F05d (.D(1'b0),.RN(frontend_0_n_91),.CK(frontend_0_n_21),.Q(inst_ad[5]),.QN());
	DFFR_X1_LVT frontend_0inst_ad_reg___05F05b3___05F05d (.D(1'b0),.RN(frontend_0_n_91),.CK(frontend_0_n_21),.Q(inst_ad[3]),.QN());
	DFFR_X1_LVT frontend_0inst_ad_reg___05F05b2___05F05d (.D(1'b0),.RN(frontend_0_n_91),.CK(frontend_0_n_21),.Q(inst_ad[2]),.QN());
	DFFR_X1_LVT frontend_0inst_ad_reg___05F05b0___05F05d (.D(frontend_0_n_18),.RN(frontend_0_n_91),.CK(frontend_0_n_21),.Q(inst_ad[0]),.QN());
	INV_X1_LVT frontend_0i_12_0 (.A(frontend_0_inst_type_nxt),.ZN(frontend_0_n_12_0));
	NAND2_X1_LVT frontend_0i_12_23 (.A1(frontend_0_n_12_8),.A2(frontend_0_n_12_0),.ZN(frontend_0_n_12_14));
	NAND3_X1_LVT frontend_0i_12_5 (.A1(frontend_0_n_12_2),.A2(frontend_0_n_12_3),.A3(frontend_0_n_12_4),.ZN(frontend_0_n_12_5));
	NOR2_X1_LVT frontend_0i_12_24 (.A1(frontend_0_n_12_14),.A2(frontend_0_n_12_5),.ZN(frontend_0_inst_as_nxt[9]));
	NOR2_X1_LVT frontend_0i_12_25 (.A1(frontend_0_n_12_14),.A2(frontend_0_n_12_3),.ZN(frontend_0_inst_as_nxt[10]));
	NOR2_X1_LVT frontend_0i_12_26 (.A1(frontend_0_n_12_14),.A2(frontend_0_n_12_2),.ZN(frontend_0_inst_as_nxt[11]));
	NOR2_X1_LVT frontend_0i_12_27 (.A1(frontend_0_n_12_14),.A2(frontend_0_n_12_4),.ZN(frontend_0_inst_as_nxt[12]));
	NOR4_X1_LVT frontend_0i_13_0 (.A1(frontend_0_inst_as_nxt[9]),.A2(frontend_0_inst_as_nxt[10]),.A3(frontend_0_inst_as_nxt[11]),.A4(frontend_0_inst_as_nxt[12]),.ZN(frontend_0_n_13_0));
	NOR3_X1_LVT frontend_0i_12_21 (.A1(frontend_0_n_12_13),.A2(frontend_0_n_12_9),.A3(frontend_0_n_12_2),.ZN(frontend_0_inst_as_nxt[7]));
	NOR3_X1_LVT frontend_0i_12_22 (.A1(frontend_0_n_12_13),.A2(frontend_0_n_12_9),.A3(frontend_0_n_12_4),.ZN(frontend_0_inst_as_nxt[8]));
	NOR2_X1_LVT frontend_0i_13_1 (.A1(frontend_0_inst_as_nxt[7]),.A2(frontend_0_inst_as_nxt[8]),.ZN(frontend_0_n_13_1));
	NAND2_X1_LVT frontend_0i_13_2 (.A1(frontend_0_n_13_0),.A2(frontend_0_n_13_1),.ZN(frontend_0_is_const));
	DFFR_X1_LVT frontend_0inst_as_reg___05F05b7___05F05d (.D(frontend_0_is_const),.RN(frontend_0_n_91),.CK(frontend_0_n_12),.Q(inst_as[7]),.QN());
	DFFR_X1_LVT frontend_0inst_as_reg___05F05b3___05F05d (.D(frontend_0_inst_as_nxt[3]),.RN(frontend_0_n_91),.CK(frontend_0_n_12),.Q(inst_as[3]),.QN());
	DFFR_X1_LVT frontend_0inst_as_reg___05F05b2___05F05d (.D(frontend_0_inst_as_nxt[2]),.RN(frontend_0_n_91),.CK(frontend_0_n_12),.Q(inst_as[2]),.QN());
	OAI21_X1_LVT frontend_0i_12_10 (.A(frontend_0_n_12_0),.B1(frontend_0_n_12_5),.B2(frontend_0_n_12_9),.ZN(frontend_0_inst_as_nxt[0]));
	DFFR_X1_LVT frontend_0inst_as_reg___05F05b0___05F05d (.D(frontend_0_inst_as_nxt[0]),.RN(frontend_0_n_91),.CK(frontend_0_n_12),.Q(inst_as[0]),.QN());
	INV_X1_LVT frontend_0i_82_1 (.A(fe_mdb_in[13]),.ZN(frontend_0_n_82_1));
	NAND2_X1_LVT frontend_0i_82_3 (.A1(fe_mdb_in[12]),.A2(frontend_0_n_82_1),.ZN(frontend_0_n_82_3));
	INV_X1_LVT frontend_0i_82_6 (.A(fe_mdb_in[14]),.ZN(frontend_0_n_82_6));
	NAND2_X1_LVT frontend_0i_82_9 (.A1(frontend_0_n_82_6),.A2(fe_mdb_in[15]),.ZN(frontend_0_n_82_9));
	NOR2_X1_LVT frontend_0i_82_16 (.A1(frontend_0_n_82_3),.A2(frontend_0_n_82_9),.ZN(frontend_0_n_98));
	AND2_X1_LVT frontend_0i_83_5 (.A1(frontend_0_n_17),.A2(frontend_0_n_98),.ZN(frontend_0_inst_to_nxt[5]));
	NAND2_X1_LVT frontend_0i_82_5 (.A1(fe_mdb_in[12]),.A2(fe_mdb_in[13]),.ZN(frontend_0_n_82_5));
	NOR2_X1_LVT frontend_0i_82_18 (.A1(frontend_0_n_82_5),.A2(frontend_0_n_82_9),.ZN(frontend_0_n_100));
	AND2_X1_LVT frontend_0i_83_7 (.A1(frontend_0_n_17),.A2(frontend_0_n_100),.ZN(frontend_0_inst_to_nxt[7]));
	OR2_X1_LVT frontend_0i_88_9 (.A1(frontend_0_inst_to_nxt[5]),.A2(frontend_0_inst_to_nxt[7]),.ZN(frontend_0_inst_alu_nxt[11]));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_alu_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_108));
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b11___05F05d (.D(frontend_0_inst_alu_nxt[11]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[11]),.QN());
	NOR2_X1_LVT frontend_0i_25_9 (.A1(frontend_0_n_25_4),.A2(fe_mdb_in[9]),.ZN(frontend_0_n_24));
	AND2_X1_LVT frontend_0i_26_2 (.A1(frontend_0_n_10),.A2(frontend_0_n_24),.ZN(frontend_0_n_32));
	AND2_X1_LVT frontend_0i_27_3 (.A1(frontend_0_n_27_0),.A2(frontend_0_n_32),.ZN(frontend_0_inst_so_nxt[2]));
	NOR2_X1_LVT frontend_0i_25_7 (.A1(frontend_0_n_25_2),.A2(fe_mdb_in[9]),.ZN(frontend_0_n_22));
	AND2_X1_LVT frontend_0i_26_0 (.A1(frontend_0_n_22),.A2(frontend_0_n_10),.ZN(frontend_0_n_30));
	AND2_X1_LVT frontend_0i_27_1 (.A1(frontend_0_n_27_0),.A2(frontend_0_n_30),.ZN(frontend_0_inst_so_nxt[0]));
	NOR2_X1_LVT frontend_0i_88_6 (.A1(frontend_0_inst_so_nxt[2]),.A2(frontend_0_inst_so_nxt[0]),.ZN(frontend_0_n_88_1));
	INV_X1_LVT frontend_0i_88_8 (.A(frontend_0_n_88_1),.ZN(frontend_0_inst_alu_nxt[10]));
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b10___05F05d (.D(frontend_0_inst_alu_nxt[10]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[10]),.QN());
	NAND2_X1_LVT frontend_0i_82_10 (.A1(fe_mdb_in[14]),.A2(fe_mdb_in[15]),.ZN(frontend_0_n_82_10));
	NOR2_X1_LVT frontend_0i_82_22 (.A1(frontend_0_n_82_5),.A2(frontend_0_n_82_10),.ZN(frontend_0_n_104));
	AND2_X1_LVT frontend_0i_83_11 (.A1(frontend_0_n_17),.A2(frontend_0_n_104),.ZN(frontend_0_inst_to_nxt[11]));
	OR2_X1_LVT frontend_0i_87_0 (.A1(frontend_0_inst_to_nxt[7]),.A2(frontend_0_inst_to_nxt[11]),.ZN(frontend_0_n_107));
	NOR2_X1_LVT frontend_0i_25_10 (.A1(frontend_0_n_25_5),.A2(fe_mdb_in[9]),.ZN(frontend_0_n_25));
	AND2_X1_LVT frontend_0i_26_3 (.A1(frontend_0_n_10),.A2(frontend_0_n_25),.ZN(frontend_0_n_33));
	AND2_X1_LVT frontend_0i_27_4 (.A1(frontend_0_n_27_0),.A2(frontend_0_n_33),.ZN(frontend_0_inst_so_nxt[3]));
	OR2_X1_LVT frontend_0i_88_4 (.A1(frontend_0_n_107),.A2(frontend_0_inst_so_nxt[3]),.ZN(frontend_0_inst_alu_nxt[8]));
	INV_X1_LVT frontend_0i_82_7 (.A(fe_mdb_in[15]),.ZN(frontend_0_n_82_7));
	NAND2_X1_LVT frontend_0i_82_8 (.A1(fe_mdb_in[14]),.A2(frontend_0_n_82_7),.ZN(frontend_0_n_82_8));
	NOR2_X1_LVT frontend_0i_82_12 (.A1(frontend_0_n_82_3),.A2(frontend_0_n_82_8),.ZN(frontend_0_n_94));
	AND2_X1_LVT frontend_0i_83_1 (.A1(frontend_0_n_17),.A2(frontend_0_n_94),.ZN(frontend_0_inst_to_nxt[1]));
	INV_X1_LVT frontend_0i_82_0 (.A(fe_mdb_in[12]),.ZN(frontend_0_n_82_0));
	NAND2_X1_LVT frontend_0i_82_2 (.A1(frontend_0_n_82_0),.A2(frontend_0_n_82_1),.ZN(frontend_0_n_82_2));
	NOR2_X1_LVT frontend_0i_82_15 (.A1(frontend_0_n_82_2),.A2(frontend_0_n_82_9),.ZN(frontend_0_n_97));
	AND2_X1_LVT frontend_0i_83_4 (.A1(frontend_0_n_17),.A2(frontend_0_n_97),.ZN(frontend_0_inst_to_nxt[4]));
	OR2_X1_LVT frontend_0i_84_0 (.A1(frontend_0_inst_to_nxt[5]),.A2(frontend_0_inst_to_nxt[4]),.ZN(frontend_0_alu_inc));
	NOR2_X1_LVT frontend_0i_82_14 (.A1(frontend_0_n_82_5),.A2(frontend_0_n_82_8),.ZN(frontend_0_n_96));
	AND2_X1_LVT frontend_0i_83_3 (.A1(frontend_0_n_17),.A2(frontend_0_n_96),.ZN(frontend_0_inst_to_nxt[3]));
	NAND2_X1_LVT frontend_0i_82_4 (.A1(frontend_0_n_82_0),.A2(fe_mdb_in[13]),.ZN(frontend_0_n_82_4));
	NOR2_X1_LVT frontend_0i_82_13 (.A1(frontend_0_n_82_4),.A2(frontend_0_n_82_8),.ZN(frontend_0_n_95));
	AND2_X1_LVT frontend_0i_83_2 (.A1(frontend_0_n_17),.A2(frontend_0_n_95),.ZN(frontend_0_inst_to_nxt[2]));
	OR2_X1_LVT frontend_0i_85_0 (.A1(frontend_0_inst_to_nxt[3]),.A2(frontend_0_inst_to_nxt[2]),.ZN(frontend_0_n_105));
	OR3_X1_LVT frontend_0i_86_0 (.A1(frontend_0_inst_to_nxt[1]),.A2(frontend_0_alu_inc),.A3(frontend_0_n_105),.ZN(frontend_0_n_106));
	NOR2_X1_LVT frontend_0i_82_21 (.A1(frontend_0_n_82_4),.A2(frontend_0_n_82_10),.ZN(frontend_0_n_103));
	AND2_X1_LVT frontend_0i_83_10 (.A1(frontend_0_n_17),.A2(frontend_0_n_103),.ZN(frontend_0_inst_to_nxt[10]));
	NOR2_X1_LVT frontend_0i_82_17 (.A1(frontend_0_n_82_4),.A2(frontend_0_n_82_9),.ZN(frontend_0_n_99));
	AND2_X1_LVT frontend_0i_83_6 (.A1(frontend_0_n_17),.A2(frontend_0_n_99),.ZN(frontend_0_inst_to_nxt[6]));
	NOR4_X1_LVT frontend_0i_88_5 (.A1(frontend_0_inst_alu_nxt[8]),.A2(frontend_0_n_106),.A3(frontend_0_inst_to_nxt[10]),.A4(frontend_0_inst_to_nxt[6]),.ZN(frontend_0_n_88_0));
	NAND2_X1_LVT frontend_0i_88_7 (.A1(frontend_0_n_88_0),.A2(frontend_0_n_88_1),.ZN(frontend_0_inst_alu_nxt[9]));
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b9___05F05d (.D(frontend_0_inst_alu_nxt[9]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[9]),.QN());
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b8___05F05d (.D(frontend_0_inst_alu_nxt[8]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[8]),.QN());
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b7___05F05d (.D(frontend_0_inst_to_nxt[6]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[7]),.QN());
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b6___05F05d (.D(frontend_0_inst_to_nxt[10]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[6]),.QN());
	NOR2_X1_LVT frontend_0i_82_20 (.A1(frontend_0_n_82_3),.A2(frontend_0_n_82_10),.ZN(frontend_0_n_102));
	AND2_X1_LVT frontend_0i_83_9 (.A1(frontend_0_n_17),.A2(frontend_0_n_102),.ZN(frontend_0_inst_to_nxt[9]));
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b5___05F05d (.D(frontend_0_inst_to_nxt[9]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[5]),.QN());
	NOR2_X1_LVT frontend_0i_82_19 (.A1(frontend_0_n_82_2),.A2(frontend_0_n_82_10),.ZN(frontend_0_n_101));
	AND2_X1_LVT frontend_0i_83_8 (.A1(frontend_0_n_17),.A2(frontend_0_n_101),.ZN(frontend_0_inst_to_nxt[8]));
	OR2_X1_LVT frontend_0i_88_3 (.A1(frontend_0_inst_to_nxt[8]),.A2(frontend_0_n_107),.ZN(frontend_0_inst_alu_nxt[4]));
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b4___05F05d (.D(frontend_0_inst_alu_nxt[4]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[4]),.QN());
	OR2_X1_LVT frontend_0i_88_2 (.A1(frontend_0_n_49),.A2(frontend_0_n_106),.ZN(frontend_0_inst_alu_nxt[3]));
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b3___05F05d (.D(frontend_0_inst_alu_nxt[3]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[3]),.QN());
	OR2_X1_LVT frontend_0i_88_1 (.A1(frontend_0_inst_to_nxt[6]),.A2(frontend_0_n_105),.ZN(frontend_0_inst_alu_nxt[2]));
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b2___05F05d (.D(frontend_0_inst_alu_nxt[2]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[2]),.QN());
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b1___05F05d (.D(frontend_0_alu_inc),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[1]),.QN());
	OR3_X1_LVT frontend_0i_88_0 (.A1(frontend_0_inst_to_nxt[3]),.A2(frontend_0_alu_inc),.A3(frontend_0_inst_to_nxt[8]),.ZN(frontend_0_inst_alu_nxt[0]));
	DFFR_X1_LVT frontend_0inst_alu_reg___05F05b0___05F05d (.D(frontend_0_inst_alu_nxt[0]),.RN(frontend_0_n_91),.CK(frontend_0_n_108),.Q(inst_alu[0]),.QN());
	NAND3_X1_LVT frontend_0i_91_0 (.A1(fe_mdb_in[6]),.A2(frontend_0_n_0),.A3(frontend_0_n_9),.ZN(frontend_0_n_91_0));
	NOR2_X1_LVT frontend_0i_91_1 (.A1(frontend_0_n_91_0),.A2(frontend_0_inst_type_nxt),.ZN(frontend_0_n_110));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_bw_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_109));
	DFFR_X1_LVT frontend_0inst_bw_reg (.D(frontend_0_n_110),.RN(frontend_0_n_91),.CK(frontend_0_n_109),.Q(inst_bw),.QN());
	DFFR_X1_LVT frontend_0inst_type_reg___05F05b1___05F05d (.D(frontend_0_inst_type_nxt),.RN(frontend_0_n_91),.CK(frontend_0_n_43),.Q(inst_type[1]),.QN());
	NOR2_X1_LVT frontend_0i_97_0 (.A1(inst_type[1]),.A2(cpu_halt_st),.ZN(frontend_0_n_97_0));
	INV_X1_LVT frontend_0i_97_1 (.A(frontend_0_n_97_0),.ZN(frontend_0_n_97_1));
	DFFR_X1_LVT frontend_0inst_so_reg___05F05b7___05F05d (.D(frontend_0_inst_so_nxt[7]),.RN(frontend_0_n_91),.CK(frontend_0_n_38),.Q(inst_so[7]),.QN());
	OR2_X1_LVT frontend_0i_96_0 (.A1(inst_so[7]),.A2(frontend_0_n_39),.ZN(frontend_0_n_144));
	NOR2_X1_LVT frontend_0i_97_2 (.A1(frontend_0_n_97_1),.A2(frontend_0_n_144),.ZN(frontend_0_n_97_2));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_dest_bin_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_111));
	DFFR_X1_LVT frontend_0inst_dest_bin_reg___05F05b0___05F05d (.D(fe_mdb_in[0]),.RN(frontend_0_n_91),.CK(frontend_0_n_111),.Q(frontend_0_inst_dest_bin[0]),.QN());
	DFFR_X1_LVT frontend_0inst_dest_bin_reg___05F05b1___05F05d (.D(fe_mdb_in[1]),.RN(frontend_0_n_91),.CK(frontend_0_n_111),.Q(frontend_0_inst_dest_bin[1]),.QN());
	NAND2_X1_LVT frontend_0i_94_5 (.A1(frontend_0_inst_dest_bin[0]),.A2(frontend_0_inst_dest_bin[1]),.ZN(frontend_0_n_94_5));
	DFFR_X1_LVT frontend_0inst_dest_bin_reg___05F05b2___05F05d (.D(fe_mdb_in[2]),.RN(frontend_0_n_91),.CK(frontend_0_n_111),.Q(frontend_0_inst_dest_bin[2]),.QN());
	DFFR_X1_LVT frontend_0inst_dest_bin_reg___05F05b3___05F05d (.D(fe_mdb_in[3]),.RN(frontend_0_n_91),.CK(frontend_0_n_111),.Q(frontend_0_inst_dest_bin[3]),.QN());
	NAND2_X1_LVT frontend_0i_94_11 (.A1(frontend_0_inst_dest_bin[2]),.A2(frontend_0_inst_dest_bin[3]),.ZN(frontend_0_n_94_11));
	NOR2_X1_LVT frontend_0i_94_27 (.A1(frontend_0_n_94_5),.A2(frontend_0_n_94_11),.ZN(frontend_0_n_127));
	NAND2_X1_LVT frontend_0i_95_5 (.A1(dbg_mem_addr[0]),.A2(dbg_mem_addr[1]),.ZN(frontend_0_n_95_5));
	NAND2_X1_LVT frontend_0i_95_11 (.A1(dbg_mem_addr[2]),.A2(dbg_mem_addr[3]),.ZN(frontend_0_n_95_11));
	NOR2_X1_LVT frontend_0i_95_27 (.A1(frontend_0_n_95_5),.A2(frontend_0_n_95_11),.ZN(frontend_0_n_143));
	AOI22_X1_LVT frontend_0i_97_34 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_127),.B1(cpu_halt_st),.B2(frontend_0_n_143),.ZN(frontend_0_n_97_19));
	INV_X1_LVT frontend_0i_97_35 (.A(frontend_0_n_97_19),.ZN(inst_dest[15]));
	INV_X1_LVT frontend_0i_94_0 (.A(frontend_0_inst_dest_bin[0]),.ZN(frontend_0_n_94_0));
	NAND2_X1_LVT frontend_0i_94_4 (.A1(frontend_0_n_94_0),.A2(frontend_0_inst_dest_bin[1]),.ZN(frontend_0_n_94_4));
	NOR2_X1_LVT frontend_0i_94_26 (.A1(frontend_0_n_94_4),.A2(frontend_0_n_94_11),.ZN(frontend_0_n_126));
	INV_X1_LVT frontend_0i_95_0 (.A(dbg_mem_addr[0]),.ZN(frontend_0_n_95_0));
	NAND2_X1_LVT frontend_0i_95_4 (.A1(frontend_0_n_95_0),.A2(dbg_mem_addr[1]),.ZN(frontend_0_n_95_4));
	NOR2_X1_LVT frontend_0i_95_26 (.A1(frontend_0_n_95_4),.A2(frontend_0_n_95_11),.ZN(frontend_0_n_142));
	AOI22_X1_LVT frontend_0i_97_32 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_126),.B1(cpu_halt_st),.B2(frontend_0_n_142),.ZN(frontend_0_n_97_18));
	INV_X1_LVT frontend_0i_97_33 (.A(frontend_0_n_97_18),.ZN(inst_dest[14]));
	INV_X1_LVT frontend_0i_94_1 (.A(frontend_0_inst_dest_bin[1]),.ZN(frontend_0_n_94_1));
	NAND2_X1_LVT frontend_0i_94_3 (.A1(frontend_0_inst_dest_bin[0]),.A2(frontend_0_n_94_1),.ZN(frontend_0_n_94_3));
	NOR2_X1_LVT frontend_0i_94_25 (.A1(frontend_0_n_94_3),.A2(frontend_0_n_94_11),.ZN(frontend_0_n_125));
	INV_X1_LVT frontend_0i_95_1 (.A(dbg_mem_addr[1]),.ZN(frontend_0_n_95_1));
	NAND2_X1_LVT frontend_0i_95_3 (.A1(dbg_mem_addr[0]),.A2(frontend_0_n_95_1),.ZN(frontend_0_n_95_3));
	NOR2_X1_LVT frontend_0i_95_25 (.A1(frontend_0_n_95_3),.A2(frontend_0_n_95_11),.ZN(frontend_0_n_141));
	AOI22_X1_LVT frontend_0i_97_30 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_125),.B1(cpu_halt_st),.B2(frontend_0_n_141),.ZN(frontend_0_n_97_17));
	INV_X1_LVT frontend_0i_97_31 (.A(frontend_0_n_97_17),.ZN(inst_dest[13]));
	NAND2_X1_LVT frontend_0i_94_2 (.A1(frontend_0_n_94_0),.A2(frontend_0_n_94_1),.ZN(frontend_0_n_94_2));
	NOR2_X1_LVT frontend_0i_94_24 (.A1(frontend_0_n_94_2),.A2(frontend_0_n_94_11),.ZN(frontend_0_n_124));
	NAND2_X1_LVT frontend_0i_95_2 (.A1(frontend_0_n_95_0),.A2(frontend_0_n_95_1),.ZN(frontend_0_n_95_2));
	NOR2_X1_LVT frontend_0i_95_24 (.A1(frontend_0_n_95_2),.A2(frontend_0_n_95_11),.ZN(frontend_0_n_140));
	AOI22_X1_LVT frontend_0i_97_28 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_124),.B1(cpu_halt_st),.B2(frontend_0_n_140),.ZN(frontend_0_n_97_16));
	INV_X1_LVT frontend_0i_97_29 (.A(frontend_0_n_97_16),.ZN(inst_dest[12]));
	INV_X1_LVT frontend_0i_94_6 (.A(frontend_0_inst_dest_bin[2]),.ZN(frontend_0_n_94_6));
	NAND2_X1_LVT frontend_0i_94_10 (.A1(frontend_0_n_94_6),.A2(frontend_0_inst_dest_bin[3]),.ZN(frontend_0_n_94_10));
	NOR2_X1_LVT frontend_0i_94_23 (.A1(frontend_0_n_94_5),.A2(frontend_0_n_94_10),.ZN(frontend_0_n_123));
	INV_X1_LVT frontend_0i_95_6 (.A(dbg_mem_addr[2]),.ZN(frontend_0_n_95_6));
	NAND2_X1_LVT frontend_0i_95_10 (.A1(frontend_0_n_95_6),.A2(dbg_mem_addr[3]),.ZN(frontend_0_n_95_10));
	NOR2_X1_LVT frontend_0i_95_23 (.A1(frontend_0_n_95_5),.A2(frontend_0_n_95_10),.ZN(frontend_0_n_139));
	AOI22_X1_LVT frontend_0i_97_26 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_123),.B1(cpu_halt_st),.B2(frontend_0_n_139),.ZN(frontend_0_n_97_15));
	INV_X1_LVT frontend_0i_97_27 (.A(frontend_0_n_97_15),.ZN(inst_dest[11]));
	NOR2_X1_LVT frontend_0i_94_22 (.A1(frontend_0_n_94_4),.A2(frontend_0_n_94_10),.ZN(frontend_0_n_122));
	NOR2_X1_LVT frontend_0i_95_22 (.A1(frontend_0_n_95_4),.A2(frontend_0_n_95_10),.ZN(frontend_0_n_138));
	AOI22_X1_LVT frontend_0i_97_24 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_122),.B1(cpu_halt_st),.B2(frontend_0_n_138),.ZN(frontend_0_n_97_14));
	INV_X1_LVT frontend_0i_97_25 (.A(frontend_0_n_97_14),.ZN(inst_dest[10]));
	NOR2_X1_LVT frontend_0i_94_21 (.A1(frontend_0_n_94_3),.A2(frontend_0_n_94_10),.ZN(frontend_0_n_121));
	NOR2_X1_LVT frontend_0i_95_21 (.A1(frontend_0_n_95_3),.A2(frontend_0_n_95_10),.ZN(frontend_0_n_137));
	AOI22_X1_LVT frontend_0i_97_22 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_121),.B1(cpu_halt_st),.B2(frontend_0_n_137),.ZN(frontend_0_n_97_13));
	INV_X1_LVT frontend_0i_97_23 (.A(frontend_0_n_97_13),.ZN(inst_dest[9]));
	NOR2_X1_LVT frontend_0i_94_20 (.A1(frontend_0_n_94_2),.A2(frontend_0_n_94_10),.ZN(frontend_0_n_120));
	NOR2_X1_LVT frontend_0i_95_20 (.A1(frontend_0_n_95_2),.A2(frontend_0_n_95_10),.ZN(frontend_0_n_136));
	AOI22_X1_LVT frontend_0i_97_20 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_120),.B1(cpu_halt_st),.B2(frontend_0_n_136),.ZN(frontend_0_n_97_12));
	INV_X1_LVT frontend_0i_97_21 (.A(frontend_0_n_97_12),.ZN(inst_dest[8]));
	INV_X1_LVT frontend_0i_94_7 (.A(frontend_0_inst_dest_bin[3]),.ZN(frontend_0_n_94_7));
	NAND2_X1_LVT frontend_0i_94_9 (.A1(frontend_0_inst_dest_bin[2]),.A2(frontend_0_n_94_7),.ZN(frontend_0_n_94_9));
	NOR2_X1_LVT frontend_0i_94_19 (.A1(frontend_0_n_94_5),.A2(frontend_0_n_94_9),.ZN(frontend_0_n_119));
	INV_X1_LVT frontend_0i_95_7 (.A(dbg_mem_addr[3]),.ZN(frontend_0_n_95_7));
	NAND2_X1_LVT frontend_0i_95_9 (.A1(dbg_mem_addr[2]),.A2(frontend_0_n_95_7),.ZN(frontend_0_n_95_9));
	NOR2_X1_LVT frontend_0i_95_19 (.A1(frontend_0_n_95_5),.A2(frontend_0_n_95_9),.ZN(frontend_0_n_135));
	AOI22_X1_LVT frontend_0i_97_18 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_119),.B1(cpu_halt_st),.B2(frontend_0_n_135),.ZN(frontend_0_n_97_11));
	INV_X1_LVT frontend_0i_97_19 (.A(frontend_0_n_97_11),.ZN(inst_dest[7]));
	NOR2_X1_LVT frontend_0i_94_18 (.A1(frontend_0_n_94_4),.A2(frontend_0_n_94_9),.ZN(frontend_0_n_118));
	NOR2_X1_LVT frontend_0i_95_18 (.A1(frontend_0_n_95_4),.A2(frontend_0_n_95_9),.ZN(frontend_0_n_134));
	AOI22_X1_LVT frontend_0i_97_16 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_118),.B1(cpu_halt_st),.B2(frontend_0_n_134),.ZN(frontend_0_n_97_10));
	INV_X1_LVT frontend_0i_97_17 (.A(frontend_0_n_97_10),.ZN(inst_dest[6]));
	NOR2_X1_LVT frontend_0i_94_17 (.A1(frontend_0_n_94_3),.A2(frontend_0_n_94_9),.ZN(frontend_0_n_117));
	NOR2_X1_LVT frontend_0i_95_17 (.A1(frontend_0_n_95_3),.A2(frontend_0_n_95_9),.ZN(frontend_0_n_133));
	AOI22_X1_LVT frontend_0i_97_14 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_117),.B1(cpu_halt_st),.B2(frontend_0_n_133),.ZN(frontend_0_n_97_9));
	INV_X1_LVT frontend_0i_97_15 (.A(frontend_0_n_97_9),.ZN(inst_dest[5]));
	NOR2_X1_LVT frontend_0i_94_16 (.A1(frontend_0_n_94_2),.A2(frontend_0_n_94_9),.ZN(frontend_0_n_116));
	NOR2_X1_LVT frontend_0i_95_16 (.A1(frontend_0_n_95_2),.A2(frontend_0_n_95_9),.ZN(frontend_0_n_132));
	AOI22_X1_LVT frontend_0i_97_12 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_116),.B1(cpu_halt_st),.B2(frontend_0_n_132),.ZN(frontend_0_n_97_8));
	INV_X1_LVT frontend_0i_97_13 (.A(frontend_0_n_97_8),.ZN(inst_dest[4]));
	NAND2_X1_LVT frontend_0i_94_8 (.A1(frontend_0_n_94_6),.A2(frontend_0_n_94_7),.ZN(frontend_0_n_94_8));
	NOR2_X1_LVT frontend_0i_94_15 (.A1(frontend_0_n_94_5),.A2(frontend_0_n_94_8),.ZN(frontend_0_n_115));
	NAND2_X1_LVT frontend_0i_95_8 (.A1(frontend_0_n_95_6),.A2(frontend_0_n_95_7),.ZN(frontend_0_n_95_8));
	NOR2_X1_LVT frontend_0i_95_15 (.A1(frontend_0_n_95_5),.A2(frontend_0_n_95_8),.ZN(frontend_0_n_131));
	AOI22_X1_LVT frontend_0i_97_10 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_115),.B1(cpu_halt_st),.B2(frontend_0_n_131),.ZN(frontend_0_n_97_7));
	INV_X1_LVT frontend_0i_97_11 (.A(frontend_0_n_97_7),.ZN(inst_dest[3]));
	NOR2_X1_LVT frontend_0i_94_14 (.A1(frontend_0_n_94_4),.A2(frontend_0_n_94_8),.ZN(frontend_0_n_114));
	NOR2_X1_LVT frontend_0i_95_14 (.A1(frontend_0_n_95_4),.A2(frontend_0_n_95_8),.ZN(frontend_0_n_130));
	AOI22_X1_LVT frontend_0i_97_8 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_114),.B1(cpu_halt_st),.B2(frontend_0_n_130),.ZN(frontend_0_n_97_6));
	INV_X1_LVT frontend_0i_97_9 (.A(frontend_0_n_97_6),.ZN(inst_dest[2]));
	NOR2_X1_LVT frontend_0i_94_13 (.A1(frontend_0_n_94_3),.A2(frontend_0_n_94_8),.ZN(frontend_0_n_113));
	NOR2_X1_LVT frontend_0i_95_13 (.A1(frontend_0_n_95_3),.A2(frontend_0_n_95_8),.ZN(frontend_0_n_129));
	AOI222_X1_LVT frontend_0i_97_6 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_113),.B1(frontend_0_n_97_0),.B2(frontend_0_n_144),.C1(cpu_halt_st),.C2(frontend_0_n_129),.ZN(frontend_0_n_97_5));
	INV_X1_LVT frontend_0i_97_7 (.A(frontend_0_n_97_5),.ZN(inst_dest[1]));
	NOR2_X1_LVT frontend_0i_94_12 (.A1(frontend_0_n_94_2),.A2(frontend_0_n_94_8),.ZN(frontend_0_n_112));
	INV_X1_LVT frontend_0i_97_3 (.A(cpu_halt_st),.ZN(frontend_0_n_97_3));
	NOR2_X1_LVT frontend_0i_95_12 (.A1(frontend_0_n_95_2),.A2(frontend_0_n_95_8),.ZN(frontend_0_n_128));
	AOI222_X1_LVT frontend_0i_97_4 (.A1(frontend_0_n_97_2),.A2(frontend_0_n_112),.B1(frontend_0_n_97_3),.B2(inst_type[1]),.C1(frontend_0_n_128),.C2(cpu_halt_st),.ZN(frontend_0_n_97_4));
	INV_X1_LVT frontend_0i_97_5 (.A(frontend_0_n_97_4),.ZN(inst_dest[0]));
	INV_X1_LVT frontend_0i_99_6 (.A(fe_mdb_in[3]),.ZN(frontend_0_n_99_4));
	XNOR2_X1_LVT frontend_0i_99_19 (.A(fe_mdb_in[15]),.B(frontend_0_n_99_4),.ZN(frontend_0_n_99_17));
	INV_X1_LVT frontend_0i_98_0 (.A(frontend_0_i_state_nxt_reg[2]),.ZN(frontend_0_n_98_0));
	OR3_X1_LVT frontend_0i_98_1 (.A1(frontend_0_n_98_0),.A2(frontend_0_i_state_nxt_reg[0]),.A3(frontend_0_i_state_nxt_reg[1]),.ZN(frontend_0_n_98_1));
	INV_X1_LVT frontend_0i_98_2 (.A(inst_as[4]),.ZN(frontend_0_n_98_2));
	AND4_X1_LVT frontend_0i_98_3 (.A1(frontend_0_n_98_1),.A2(frontend_0_n_98_2),.A3(frontend_0_n_6),.A4(inst_ad[4]),.ZN(frontend_0_n_98_3));
	AOI221_X1_LVT frontend_0i_98_4 (.A(frontend_0_n_98_3),.B1(frontend_0_n_6),.B2(inst_as[4]),.C1(frontend_0_n_7),.C2(inst_ad[4]),.ZN(frontend_0_n_98_4));
	INV_X1_LVT frontend_0i_98_5 (.A(frontend_0_n_98_4),.ZN(frontend_0_n_145));
	INV_X1_LVT frontend_0i_99_3 (.A(fe_mdb_in[1]),.ZN(frontend_0_n_99_2));
	NAND2_X1_LVT frontend_0i_99_2 (.A1(frontend_0_n_145),.A2(frontend_0_n_99_2),.ZN(frontend_0_n_99_1));
	OR2_X1_LVT frontend_0i_99_5 (.A1(fe_mdb_in[2]),.A2(frontend_0_n_99_1),.ZN(frontend_0_n_99_3));
	HA_X1_LVT frontend_0i_99_7 (.A(frontend_0_n_99_4),.B(frontend_0_n_99_3),.CO(frontend_0_n_99_5),.S(frontend_0_ext_nxt[3]));
	FA_X1_LVT frontend_0i_99_8 (.A(fe_mdb_in[4]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_5),.CO(frontend_0_n_99_6),.S(frontend_0_ext_nxt[4]));
	FA_X1_LVT frontend_0i_99_9 (.A(fe_mdb_in[5]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_6),.CO(frontend_0_n_99_7),.S(frontend_0_ext_nxt[5]));
	FA_X1_LVT frontend_0i_99_10 (.A(fe_mdb_in[6]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_7),.CO(frontend_0_n_99_8),.S(frontend_0_ext_nxt[6]));
	FA_X1_LVT frontend_0i_99_11 (.A(fe_mdb_in[7]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_8),.CO(frontend_0_n_99_9),.S(frontend_0_ext_nxt[7]));
	FA_X1_LVT frontend_0i_99_12 (.A(fe_mdb_in[8]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_9),.CO(frontend_0_n_99_10),.S(frontend_0_ext_nxt[8]));
	FA_X1_LVT frontend_0i_99_13 (.A(fe_mdb_in[9]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_10),.CO(frontend_0_n_99_11),.S(frontend_0_ext_nxt[9]));
	FA_X1_LVT frontend_0i_99_14 (.A(fe_mdb_in[10]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_11),.CO(frontend_0_n_99_12),.S(frontend_0_ext_nxt[10]));
	FA_X1_LVT frontend_0i_99_15 (.A(fe_mdb_in[11]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_12),.CO(frontend_0_n_99_13),.S(frontend_0_ext_nxt[11]));
	FA_X1_LVT frontend_0i_99_16 (.A(fe_mdb_in[12]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_13),.CO(frontend_0_n_99_14),.S(frontend_0_ext_nxt[12]));
	FA_X1_LVT frontend_0i_99_17 (.A(fe_mdb_in[13]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_14),.CO(frontend_0_n_99_15),.S(frontend_0_ext_nxt[13]));
	FA_X1_LVT frontend_0i_99_18 (.A(fe_mdb_in[14]),.B(frontend_0_n_99_4),.CI(frontend_0_n_99_15),.CO(frontend_0_n_99_16),.S(frontend_0_ext_nxt[14]));
	XNOR2_X1_LVT frontend_0i_99_20 (.A(frontend_0_n_99_17),.B(frontend_0_n_99_16),.ZN(frontend_0_ext_nxt[15]));
	INV_X1_LVT frontend_0i_101_0 (.A(frontend_0_i_state[2]),.ZN(frontend_0_n_101_0));
	NOR3_X1_LVT frontend_0i_101_1 (.A1(frontend_0_n_101_0),.A2(frontend_0_i_state[0]),.A3(frontend_0_i_state[1]),.ZN(frontend_0_n_101_1));
	OR2_X1_LVT frontend_0i_101_2 (.A1(frontend_0_n_101_1),.A2(frontend_0_n_13),.ZN(frontend_0_n_147));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_dext_reg (.CK(cpu_mclk),.E(frontend_0_n_147),.SE(1'b0),.GCK(frontend_0_n_146));
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b15___05F05d (.D(frontend_0_ext_nxt[15]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[15]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b14___05F05d (.D(frontend_0_ext_nxt[14]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[14]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b13___05F05d (.D(frontend_0_ext_nxt[13]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[13]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b12___05F05d (.D(frontend_0_ext_nxt[12]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[12]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b11___05F05d (.D(frontend_0_ext_nxt[11]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[11]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b10___05F05d (.D(frontend_0_ext_nxt[10]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[10]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b9___05F05d (.D(frontend_0_ext_nxt[9]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[9]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b8___05F05d (.D(frontend_0_ext_nxt[8]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[8]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b7___05F05d (.D(frontend_0_ext_nxt[7]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[7]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b6___05F05d (.D(frontend_0_ext_nxt[6]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[6]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b5___05F05d (.D(frontend_0_ext_nxt[5]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[5]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b4___05F05d (.D(frontend_0_ext_nxt[4]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[4]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b3___05F05d (.D(frontend_0_ext_nxt[3]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[3]),.QN());
	XNOR2_X1_LVT frontend_0i_99_4 (.A(fe_mdb_in[2]),.B(frontend_0_n_99_1),.ZN(frontend_0_ext_nxt[2]));
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b2___05F05d (.D(frontend_0_ext_nxt[2]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[2]),.QN());
	XNOR2_X1_LVT frontend_0i_99_0 (.A(frontend_0_n_145),.B(fe_mdb_in[1]),.ZN(frontend_0_n_99_0));
	INV_X1_LVT frontend_0i_99_1 (.A(frontend_0_n_99_0),.ZN(frontend_0_ext_nxt[1]));
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b1___05F05d (.D(frontend_0_ext_nxt[1]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[1]),.QN());
	DFFR_X1_LVT frontend_0inst_dext_reg___05F05b0___05F05d (.D(fe_mdb_in[0]),.RN(frontend_0_n_91),.CK(frontend_0_n_146),.Q(inst_dext[0]),.QN());
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_irq_rst_reg (.CK(cpu_mclk),.E(exec_done),.SE(1'b0),.GCK(frontend_0_n_148));
	DFFS_X1_LVT frontend_0inst_irq_rst_reg (.D(1'b0),.SN(frontend_0_n_91),.CK(frontend_0_n_148),.Q(inst_irq_rst),.QN());
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_jmp_bin_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_149));
	DFFR_X1_LVT frontend_0inst_jmp_bin_reg___05F05b0___05F05d (.D(fe_mdb_in[10]),.RN(frontend_0_n_91),.CK(frontend_0_n_149),.Q(frontend_0_inst_jmp_bin[0]),.QN());
	DFFR_X1_LVT frontend_0inst_jmp_bin_reg___05F05b1___05F05d (.D(fe_mdb_in[11]),.RN(frontend_0_n_91),.CK(frontend_0_n_149),.Q(frontend_0_inst_jmp_bin[1]),.QN());
	NAND2_X1_LVT frontend_0i_105_5 (.A1(frontend_0_inst_jmp_bin[0]),.A2(frontend_0_inst_jmp_bin[1]),.ZN(frontend_0_n_105_5));
	DFFR_X1_LVT frontend_0inst_jmp_bin_reg___05F05b2___05F05d (.D(fe_mdb_in[12]),.RN(frontend_0_n_91),.CK(frontend_0_n_149),.Q(frontend_0_inst_jmp_bin[2]),.QN());
	INV_X1_LVT frontend_0i_105_6 (.A(frontend_0_inst_jmp_bin[2]),.ZN(frontend_0_n_105_6));
	NOR2_X1_LVT frontend_0i_105_14 (.A1(frontend_0_n_105_5),.A2(frontend_0_n_105_6),.ZN(frontend_0_n_157));
	AND2_X1_LVT frontend_0i_106_7 (.A1(inst_type[1]),.A2(frontend_0_n_157),.ZN(inst_jmp[7]));
	INV_X1_LVT frontend_0i_105_0 (.A(frontend_0_inst_jmp_bin[0]),.ZN(frontend_0_n_105_0));
	NAND2_X1_LVT frontend_0i_105_4 (.A1(frontend_0_n_105_0),.A2(frontend_0_inst_jmp_bin[1]),.ZN(frontend_0_n_105_4));
	NOR2_X1_LVT frontend_0i_105_13 (.A1(frontend_0_n_105_4),.A2(frontend_0_n_105_6),.ZN(frontend_0_n_156));
	AND2_X1_LVT frontend_0i_106_6 (.A1(inst_type[1]),.A2(frontend_0_n_156),.ZN(inst_jmp[6]));
	INV_X1_LVT frontend_0i_105_1 (.A(frontend_0_inst_jmp_bin[1]),.ZN(frontend_0_n_105_1));
	NAND2_X1_LVT frontend_0i_105_3 (.A1(frontend_0_inst_jmp_bin[0]),.A2(frontend_0_n_105_1),.ZN(frontend_0_n_105_3));
	NOR2_X1_LVT frontend_0i_105_12 (.A1(frontend_0_n_105_3),.A2(frontend_0_n_105_6),.ZN(frontend_0_n_155));
	AND2_X1_LVT frontend_0i_106_5 (.A1(inst_type[1]),.A2(frontend_0_n_155),.ZN(inst_jmp[5]));
	NAND2_X1_LVT frontend_0i_105_2 (.A1(frontend_0_n_105_0),.A2(frontend_0_n_105_1),.ZN(frontend_0_n_105_2));
	NOR2_X1_LVT frontend_0i_105_11 (.A1(frontend_0_n_105_2),.A2(frontend_0_n_105_6),.ZN(frontend_0_n_154));
	AND2_X1_LVT frontend_0i_106_4 (.A1(inst_type[1]),.A2(frontend_0_n_154),.ZN(inst_jmp[4]));
	NOR2_X1_LVT frontend_0i_105_10 (.A1(frontend_0_n_105_5),.A2(frontend_0_inst_jmp_bin[2]),.ZN(frontend_0_n_153));
	AND2_X1_LVT frontend_0i_106_3 (.A1(inst_type[1]),.A2(frontend_0_n_153),.ZN(inst_jmp[3]));
	NOR2_X1_LVT frontend_0i_105_9 (.A1(frontend_0_n_105_4),.A2(frontend_0_inst_jmp_bin[2]),.ZN(frontend_0_n_152));
	AND2_X1_LVT frontend_0i_106_2 (.A1(inst_type[1]),.A2(frontend_0_n_152),.ZN(inst_jmp[2]));
	NOR2_X1_LVT frontend_0i_105_8 (.A1(frontend_0_n_105_3),.A2(frontend_0_inst_jmp_bin[2]),.ZN(frontend_0_n_151));
	AND2_X1_LVT frontend_0i_106_1 (.A1(inst_type[1]),.A2(frontend_0_n_151),.ZN(inst_jmp[1]));
	NOR2_X1_LVT frontend_0i_105_7 (.A1(frontend_0_n_105_2),.A2(frontend_0_inst_jmp_bin[2]),.ZN(frontend_0_n_150));
	AND2_X1_LVT frontend_0i_106_0 (.A1(frontend_0_n_150),.A2(inst_type[1]),.ZN(inst_jmp[0]));
	NOR2_X1_LVT frontend_0i_82_11 (.A1(frontend_0_n_82_2),.A2(frontend_0_n_82_8),.ZN(frontend_0_n_93));
	AND2_X1_LVT frontend_0i_83_0 (.A1(frontend_0_n_17),.A2(frontend_0_n_93),.ZN(frontend_0_inst_to_nxt[0]));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_mov_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_158));
	DFFR_X1_LVT frontend_0inst_mov_reg (.D(frontend_0_inst_to_nxt[0]),.RN(frontend_0_n_91),.CK(frontend_0_n_158),.Q(inst_mov),.QN());
	AND2_X1_LVT frontend_0i_110_33 (.A1(frontend_0_inst_type_nxt),.A2(fe_mdb_in[9]),.ZN(frontend_0_n_110_23));
	AND2_X1_LVT frontend_0i_110_14 (.A1(frontend_0_is_const),.A2(frontend_0_inst_as_nxt[12]),.ZN(frontend_0_n_110_10));
	NOR2_X1_LVT frontend_0i_110_0 (.A1(frontend_0_inst_type_nxt),.A2(frontend_0_is_const),.ZN(frontend_0_n_110_0));
	AOI211_X1_LVT frontend_0i_110_49 (.A(frontend_0_n_110_23),.B(frontend_0_n_110_10),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[15]),.ZN(frontend_0_n_110_34));
	INV_X1_LVT frontend_0i_110_2 (.A(frontend_0_decode),.ZN(frontend_0_n_110_2));
	INV_X1_LVT frontend_0i_110_50 (.A(frontend_0_ext_nxt[15]),.ZN(frontend_0_n_110_35));
	OAI22_X1_LVT frontend_0i_110_51 (.A1(frontend_0_n_110_34),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_35),.ZN(frontend_0_n_179));
	NOR2_X1_LVT frontend_0i_111_0 (.A1(frontend_0_inst_type_nxt),.A2(frontend_0_is_const),.ZN(frontend_0_n_111_0));
	INV_X1_LVT frontend_0i_111_4 (.A(frontend_0_n_111_0),.ZN(frontend_0_n_111_3));
	NOR2_X1_LVT frontend_0i_111_5 (.A1(frontend_0_inst_sext_rdy),.A2(frontend_0_n_111_3),.ZN(frontend_0_n_111_4));
	INV_X1_LVT frontend_0i_111_1 (.A(frontend_0_decode),.ZN(frontend_0_n_111_1));
	INV_X1_LVT frontend_0i_111_2 (.A(frontend_0_inst_sext_rdy),.ZN(frontend_0_n_111_2));
	OAI22_X1_LVT frontend_0i_111_3 (.A1(frontend_0_n_111_4),.A2(frontend_0_n_111_1),.B1(frontend_0_decode),.B2(frontend_0_n_111_2),.ZN(frontend_0_n_180));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_sext_reg (.CK(cpu_mclk),.E(frontend_0_n_180),.SE(1'b0),.GCK(frontend_0_n_163));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b15___05F05d (.D(frontend_0_n_179),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[15]),.QN());
	AOI211_X1_LVT frontend_0i_110_46 (.A(frontend_0_n_110_23),.B(frontend_0_n_110_10),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[14]),.ZN(frontend_0_n_110_32));
	INV_X1_LVT frontend_0i_110_47 (.A(frontend_0_ext_nxt[14]),.ZN(frontend_0_n_110_33));
	OAI22_X1_LVT frontend_0i_110_48 (.A1(frontend_0_n_110_32),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_33),.ZN(frontend_0_n_178));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b14___05F05d (.D(frontend_0_n_178),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[14]),.QN());
	AOI211_X1_LVT frontend_0i_110_43 (.A(frontend_0_n_110_23),.B(frontend_0_n_110_10),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[13]),.ZN(frontend_0_n_110_30));
	INV_X1_LVT frontend_0i_110_44 (.A(frontend_0_ext_nxt[13]),.ZN(frontend_0_n_110_31));
	OAI22_X1_LVT frontend_0i_110_45 (.A1(frontend_0_n_110_30),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_31),.ZN(frontend_0_n_177));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b13___05F05d (.D(frontend_0_n_177),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[13]),.QN());
	AOI211_X1_LVT frontend_0i_110_40 (.A(frontend_0_n_110_23),.B(frontend_0_n_110_10),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[12]),.ZN(frontend_0_n_110_28));
	INV_X1_LVT frontend_0i_110_41 (.A(frontend_0_ext_nxt[12]),.ZN(frontend_0_n_110_29));
	OAI22_X1_LVT frontend_0i_110_42 (.A1(frontend_0_n_110_28),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_29),.ZN(frontend_0_n_176));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b12___05F05d (.D(frontend_0_n_176),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[12]),.QN());
	AOI211_X1_LVT frontend_0i_110_37 (.A(frontend_0_n_110_23),.B(frontend_0_n_110_10),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[11]),.ZN(frontend_0_n_110_26));
	INV_X1_LVT frontend_0i_110_38 (.A(frontend_0_ext_nxt[11]),.ZN(frontend_0_n_110_27));
	OAI22_X1_LVT frontend_0i_110_39 (.A1(frontend_0_n_110_26),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_27),.ZN(frontend_0_n_175));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b11___05F05d (.D(frontend_0_n_175),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[11]),.QN());
	AOI211_X1_LVT frontend_0i_110_34 (.A(frontend_0_n_110_23),.B(frontend_0_n_110_10),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[10]),.ZN(frontend_0_n_110_24));
	INV_X1_LVT frontend_0i_110_35 (.A(frontend_0_ext_nxt[10]),.ZN(frontend_0_n_110_25));
	OAI22_X1_LVT frontend_0i_110_36 (.A1(frontend_0_n_110_24),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_25),.ZN(frontend_0_n_174));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b10___05F05d (.D(frontend_0_n_174),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[10]),.QN());
	AOI221_X1_LVT frontend_0i_110_30 (.A(frontend_0_n_110_10),.B1(frontend_0_inst_type_nxt),.B2(fe_mdb_in[8]),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[9]),.ZN(frontend_0_n_110_21));
	INV_X1_LVT frontend_0i_110_31 (.A(frontend_0_ext_nxt[9]),.ZN(frontend_0_n_110_22));
	OAI22_X1_LVT frontend_0i_110_32 (.A1(frontend_0_n_110_21),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_22),.ZN(frontend_0_n_173));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b9___05F05d (.D(frontend_0_n_173),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[9]),.QN());
	AOI221_X1_LVT frontend_0i_110_27 (.A(frontend_0_n_110_10),.B1(frontend_0_inst_type_nxt),.B2(fe_mdb_in[7]),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[8]),.ZN(frontend_0_n_110_19));
	INV_X1_LVT frontend_0i_110_28 (.A(frontend_0_ext_nxt[8]),.ZN(frontend_0_n_110_20));
	OAI22_X1_LVT frontend_0i_110_29 (.A1(frontend_0_n_110_19),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_20),.ZN(frontend_0_n_172));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b8___05F05d (.D(frontend_0_n_172),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[8]),.QN());
	AOI221_X1_LVT frontend_0i_110_24 (.A(frontend_0_n_110_10),.B1(frontend_0_inst_type_nxt),.B2(fe_mdb_in[6]),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[7]),.ZN(frontend_0_n_110_17));
	INV_X1_LVT frontend_0i_110_25 (.A(frontend_0_ext_nxt[7]),.ZN(frontend_0_n_110_18));
	OAI22_X1_LVT frontend_0i_110_26 (.A1(frontend_0_n_110_17),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_18),.ZN(frontend_0_n_171));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b7___05F05d (.D(frontend_0_n_171),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[7]),.QN());
	AOI221_X1_LVT frontend_0i_110_21 (.A(frontend_0_n_110_10),.B1(frontend_0_inst_type_nxt),.B2(fe_mdb_in[5]),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[6]),.ZN(frontend_0_n_110_15));
	INV_X1_LVT frontend_0i_110_22 (.A(frontend_0_ext_nxt[6]),.ZN(frontend_0_n_110_16));
	OAI22_X1_LVT frontend_0i_110_23 (.A1(frontend_0_n_110_15),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_16),.ZN(frontend_0_n_170));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b6___05F05d (.D(frontend_0_n_170),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[6]),.QN());
	AOI221_X1_LVT frontend_0i_110_18 (.A(frontend_0_n_110_10),.B1(frontend_0_inst_type_nxt),.B2(fe_mdb_in[4]),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[5]),.ZN(frontend_0_n_110_13));
	INV_X1_LVT frontend_0i_110_19 (.A(frontend_0_ext_nxt[5]),.ZN(frontend_0_n_110_14));
	OAI22_X1_LVT frontend_0i_110_20 (.A1(frontend_0_n_110_13),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_14),.ZN(frontend_0_n_169));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b5___05F05d (.D(frontend_0_n_169),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[5]),.QN());
	AOI221_X1_LVT frontend_0i_110_15 (.A(frontend_0_n_110_10),.B1(frontend_0_inst_type_nxt),.B2(fe_mdb_in[3]),.C1(frontend_0_n_110_0),.C2(frontend_0_ext_nxt[4]),.ZN(frontend_0_n_110_11));
	INV_X1_LVT frontend_0i_110_16 (.A(frontend_0_ext_nxt[4]),.ZN(frontend_0_n_110_12));
	OAI22_X1_LVT frontend_0i_110_17 (.A1(frontend_0_n_110_11),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_12),.ZN(frontend_0_n_168));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b4___05F05d (.D(frontend_0_n_168),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[4]),.QN());
	OR2_X1_LVT frontend_0i_108_3 (.A1(frontend_0_inst_as_nxt[12]),.A2(frontend_0_inst_as_nxt[8]),.ZN(frontend_0_n_162));
	AOI222_X1_LVT frontend_0i_110_11 (.A1(frontend_0_n_110_0),.A2(frontend_0_ext_nxt[3]),.B1(frontend_0_is_const),.B2(frontend_0_n_162),.C1(frontend_0_inst_type_nxt),.C2(fe_mdb_in[2]),.ZN(frontend_0_n_110_8));
	INV_X1_LVT frontend_0i_110_12 (.A(frontend_0_ext_nxt[3]),.ZN(frontend_0_n_110_9));
	OAI22_X1_LVT frontend_0i_110_13 (.A1(frontend_0_n_110_8),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_9),.ZN(frontend_0_n_167));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b3___05F05d (.D(frontend_0_n_167),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[3]),.QN());
	OR2_X1_LVT frontend_0i_108_2 (.A1(frontend_0_inst_as_nxt[12]),.A2(frontend_0_inst_as_nxt[7]),.ZN(frontend_0_n_161));
	AOI222_X1_LVT frontend_0i_110_8 (.A1(frontend_0_n_110_0),.A2(frontend_0_ext_nxt[2]),.B1(frontend_0_is_const),.B2(frontend_0_n_161),.C1(frontend_0_inst_type_nxt),.C2(fe_mdb_in[1]),.ZN(frontend_0_n_110_6));
	INV_X1_LVT frontend_0i_110_9 (.A(frontend_0_ext_nxt[2]),.ZN(frontend_0_n_110_7));
	OAI22_X1_LVT frontend_0i_110_10 (.A1(frontend_0_n_110_6),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_7),.ZN(frontend_0_n_166));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b2___05F05d (.D(frontend_0_n_166),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[2]),.QN());
	OR2_X1_LVT frontend_0i_108_1 (.A1(frontend_0_inst_as_nxt[12]),.A2(frontend_0_inst_as_nxt[11]),.ZN(frontend_0_n_160));
	AOI222_X1_LVT frontend_0i_110_5 (.A1(frontend_0_n_110_0),.A2(frontend_0_ext_nxt[1]),.B1(frontend_0_is_const),.B2(frontend_0_n_160),.C1(frontend_0_inst_type_nxt),.C2(fe_mdb_in[0]),.ZN(frontend_0_n_110_4));
	INV_X1_LVT frontend_0i_110_6 (.A(frontend_0_ext_nxt[1]),.ZN(frontend_0_n_110_5));
	OAI22_X1_LVT frontend_0i_110_7 (.A1(frontend_0_n_110_4),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_5),.ZN(frontend_0_n_165));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b1___05F05d (.D(frontend_0_n_165),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[1]),.QN());
	OR2_X1_LVT frontend_0i_108_0 (.A1(frontend_0_inst_as_nxt[12]),.A2(frontend_0_inst_as_nxt[10]),.ZN(frontend_0_n_159));
	AOI22_X1_LVT frontend_0i_110_1 (.A1(frontend_0_n_110_0),.A2(fe_mdb_in[0]),.B1(frontend_0_n_159),.B2(frontend_0_is_const),.ZN(frontend_0_n_110_1));
	INV_X1_LVT frontend_0i_110_3 (.A(fe_mdb_in[0]),.ZN(frontend_0_n_110_3));
	OAI22_X1_LVT frontend_0i_110_4 (.A1(frontend_0_n_110_1),.A2(frontend_0_n_110_2),.B1(frontend_0_decode),.B2(frontend_0_n_110_3),.ZN(frontend_0_n_164));
	DFFR_X1_LVT frontend_0inst_sext_reg___05F05b0___05F05d (.D(frontend_0_n_164),.RN(frontend_0_n_91),.CK(frontend_0_n_163),.Q(inst_sext[0]),.QN());
	DFFR_X1_LVT frontend_0inst_so_reg___05F05b3___05F05d (.D(frontend_0_inst_so_nxt[3]),.RN(frontend_0_n_91),.CK(frontend_0_n_38),.Q(inst_so[3]),.QN());
	DFFR_X1_LVT frontend_0inst_so_reg___05F05b2___05F05d (.D(frontend_0_inst_so_nxt[2]),.RN(frontend_0_n_91),.CK(frontend_0_n_38),.Q(inst_so[2]),.QN());
	NOR2_X1_LVT frontend_0i_25_8 (.A1(frontend_0_n_25_3),.A2(fe_mdb_in[9]),.ZN(frontend_0_n_23));
	AND2_X1_LVT frontend_0i_26_1 (.A1(frontend_0_n_10),.A2(frontend_0_n_23),.ZN(frontend_0_n_31));
	AND2_X1_LVT frontend_0i_27_2 (.A1(frontend_0_n_27_0),.A2(frontend_0_n_31),.ZN(frontend_0_inst_so_nxt[1]));
	DFFR_X1_LVT frontend_0inst_so_reg___05F05b1___05F05d (.D(frontend_0_inst_so_nxt[1]),.RN(frontend_0_n_91),.CK(frontend_0_n_38),.Q(inst_so[1]),.QN());
	DFFR_X1_LVT frontend_0inst_so_reg___05F05b0___05F05d (.D(frontend_0_inst_so_nxt[0]),.RN(frontend_0_n_91),.CK(frontend_0_n_38),.Q(inst_so[0]),.QN());
	DFFR_X1_LVT frontend_0inst_type_reg___05F05b2___05F05d (.D(frontend_0_n_17),.RN(frontend_0_n_91),.CK(frontend_0_n_43),.Q(inst_type[2]),.QN());
	NOR2_X1_LVT frontend_0i_115_0 (.A1(inst_so[6]),.A2(inst_type[2]),.ZN(frontend_0_n_115_0));
	INV_X1_LVT frontend_0i_115_1 (.A(inst_so[7]),.ZN(frontend_0_n_115_1));
	AND3_X1_LVT frontend_0i_115_2 (.A1(frontend_0_n_115_0),.A2(frontend_0_n_115_1),.A3(inst_type[0]),.ZN(frontend_0_n_115_2));
	CLKGATETST_X1_LVT frontend_0clk_gate_inst_src_bin_reg (.CK(cpu_mclk),.E(frontend_0_decode),.SE(1'b0),.GCK(frontend_0_n_181));
	DFFR_X1_LVT frontend_0inst_src_bin_reg___05F05b0___05F05d (.D(fe_mdb_in[8]),.RN(frontend_0_n_91),.CK(frontend_0_n_181),.Q(frontend_0_inst_src_bin[0]),.QN());
	DFFR_X1_LVT frontend_0inst_src_bin_reg___05F05b1___05F05d (.D(fe_mdb_in[9]),.RN(frontend_0_n_91),.CK(frontend_0_n_181),.Q(frontend_0_inst_src_bin[1]),.QN());
	NAND2_X1_LVT frontend_0i_114_5 (.A1(frontend_0_inst_src_bin[0]),.A2(frontend_0_inst_src_bin[1]),.ZN(frontend_0_n_114_5));
	DFFR_X1_LVT frontend_0inst_src_bin_reg___05F05b2___05F05d (.D(fe_mdb_in[10]),.RN(frontend_0_n_91),.CK(frontend_0_n_181),.Q(frontend_0_inst_src_bin[2]),.QN());
	DFFR_X1_LVT frontend_0inst_src_bin_reg___05F05b3___05F05d (.D(fe_mdb_in[11]),.RN(frontend_0_n_91),.CK(frontend_0_n_181),.Q(frontend_0_inst_src_bin[3]),.QN());
	NAND2_X1_LVT frontend_0i_114_11 (.A1(frontend_0_inst_src_bin[2]),.A2(frontend_0_inst_src_bin[3]),.ZN(frontend_0_n_114_11));
	NOR2_X1_LVT frontend_0i_114_27 (.A1(frontend_0_n_114_5),.A2(frontend_0_n_114_11),.ZN(frontend_0_n_197));
	AOI22_X1_LVT frontend_0i_115_34 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_127),.B1(inst_type[2]),.B2(frontend_0_n_197),.ZN(frontend_0_n_115_19));
	INV_X1_LVT frontend_0i_115_35 (.A(frontend_0_n_115_19),.ZN(inst_src[15]));
	INV_X1_LVT frontend_0i_114_0 (.A(frontend_0_inst_src_bin[0]),.ZN(frontend_0_n_114_0));
	NAND2_X1_LVT frontend_0i_114_4 (.A1(frontend_0_n_114_0),.A2(frontend_0_inst_src_bin[1]),.ZN(frontend_0_n_114_4));
	NOR2_X1_LVT frontend_0i_114_26 (.A1(frontend_0_n_114_4),.A2(frontend_0_n_114_11),.ZN(frontend_0_n_196));
	AOI22_X1_LVT frontend_0i_115_32 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_126),.B1(inst_type[2]),.B2(frontend_0_n_196),.ZN(frontend_0_n_115_18));
	INV_X1_LVT frontend_0i_115_33 (.A(frontend_0_n_115_18),.ZN(inst_src[14]));
	INV_X1_LVT frontend_0i_114_1 (.A(frontend_0_inst_src_bin[1]),.ZN(frontend_0_n_114_1));
	NAND2_X1_LVT frontend_0i_114_3 (.A1(frontend_0_inst_src_bin[0]),.A2(frontend_0_n_114_1),.ZN(frontend_0_n_114_3));
	NOR2_X1_LVT frontend_0i_114_25 (.A1(frontend_0_n_114_3),.A2(frontend_0_n_114_11),.ZN(frontend_0_n_195));
	AOI22_X1_LVT frontend_0i_115_30 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_125),.B1(inst_type[2]),.B2(frontend_0_n_195),.ZN(frontend_0_n_115_17));
	INV_X1_LVT frontend_0i_115_31 (.A(frontend_0_n_115_17),.ZN(inst_src[13]));
	NAND2_X1_LVT frontend_0i_114_2 (.A1(frontend_0_n_114_0),.A2(frontend_0_n_114_1),.ZN(frontend_0_n_114_2));
	NOR2_X1_LVT frontend_0i_114_24 (.A1(frontend_0_n_114_2),.A2(frontend_0_n_114_11),.ZN(frontend_0_n_194));
	AOI22_X1_LVT frontend_0i_115_28 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_124),.B1(inst_type[2]),.B2(frontend_0_n_194),.ZN(frontend_0_n_115_16));
	INV_X1_LVT frontend_0i_115_29 (.A(frontend_0_n_115_16),.ZN(inst_src[12]));
	INV_X1_LVT frontend_0i_114_6 (.A(frontend_0_inst_src_bin[2]),.ZN(frontend_0_n_114_6));
	NAND2_X1_LVT frontend_0i_114_10 (.A1(frontend_0_n_114_6),.A2(frontend_0_inst_src_bin[3]),.ZN(frontend_0_n_114_10));
	NOR2_X1_LVT frontend_0i_114_23 (.A1(frontend_0_n_114_5),.A2(frontend_0_n_114_10),.ZN(frontend_0_n_193));
	AOI22_X1_LVT frontend_0i_115_26 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_123),.B1(inst_type[2]),.B2(frontend_0_n_193),.ZN(frontend_0_n_115_15));
	INV_X1_LVT frontend_0i_115_27 (.A(frontend_0_n_115_15),.ZN(inst_src[11]));
	NOR2_X1_LVT frontend_0i_114_22 (.A1(frontend_0_n_114_4),.A2(frontend_0_n_114_10),.ZN(frontend_0_n_192));
	AOI22_X1_LVT frontend_0i_115_24 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_122),.B1(inst_type[2]),.B2(frontend_0_n_192),.ZN(frontend_0_n_115_14));
	INV_X1_LVT frontend_0i_115_25 (.A(frontend_0_n_115_14),.ZN(inst_src[10]));
	NOR2_X1_LVT frontend_0i_114_21 (.A1(frontend_0_n_114_3),.A2(frontend_0_n_114_10),.ZN(frontend_0_n_191));
	AOI22_X1_LVT frontend_0i_115_22 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_121),.B1(inst_type[2]),.B2(frontend_0_n_191),.ZN(frontend_0_n_115_13));
	INV_X1_LVT frontend_0i_115_23 (.A(frontend_0_n_115_13),.ZN(inst_src[9]));
	NOR2_X1_LVT frontend_0i_114_20 (.A1(frontend_0_n_114_2),.A2(frontend_0_n_114_10),.ZN(frontend_0_n_190));
	AOI22_X1_LVT frontend_0i_115_20 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_120),.B1(inst_type[2]),.B2(frontend_0_n_190),.ZN(frontend_0_n_115_12));
	INV_X1_LVT frontend_0i_115_21 (.A(frontend_0_n_115_12),.ZN(inst_src[8]));
	INV_X1_LVT frontend_0i_114_7 (.A(frontend_0_inst_src_bin[3]),.ZN(frontend_0_n_114_7));
	NAND2_X1_LVT frontend_0i_114_9 (.A1(frontend_0_inst_src_bin[2]),.A2(frontend_0_n_114_7),.ZN(frontend_0_n_114_9));
	NOR2_X1_LVT frontend_0i_114_19 (.A1(frontend_0_n_114_5),.A2(frontend_0_n_114_9),.ZN(frontend_0_n_189));
	AOI22_X1_LVT frontend_0i_115_18 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_119),.B1(inst_type[2]),.B2(frontend_0_n_189),.ZN(frontend_0_n_115_11));
	INV_X1_LVT frontend_0i_115_19 (.A(frontend_0_n_115_11),.ZN(inst_src[7]));
	NOR2_X1_LVT frontend_0i_114_18 (.A1(frontend_0_n_114_4),.A2(frontend_0_n_114_9),.ZN(frontend_0_n_188));
	AOI22_X1_LVT frontend_0i_115_16 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_118),.B1(inst_type[2]),.B2(frontend_0_n_188),.ZN(frontend_0_n_115_10));
	INV_X1_LVT frontend_0i_115_17 (.A(frontend_0_n_115_10),.ZN(inst_src[6]));
	NOR2_X1_LVT frontend_0i_114_17 (.A1(frontend_0_n_114_3),.A2(frontend_0_n_114_9),.ZN(frontend_0_n_187));
	AOI22_X1_LVT frontend_0i_115_14 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_117),.B1(inst_type[2]),.B2(frontend_0_n_187),.ZN(frontend_0_n_115_9));
	INV_X1_LVT frontend_0i_115_15 (.A(frontend_0_n_115_9),.ZN(inst_src[5]));
	NOR2_X1_LVT frontend_0i_114_16 (.A1(frontend_0_n_114_2),.A2(frontend_0_n_114_9),.ZN(frontend_0_n_186));
	AOI22_X1_LVT frontend_0i_115_12 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_116),.B1(inst_type[2]),.B2(frontend_0_n_186),.ZN(frontend_0_n_115_8));
	INV_X1_LVT frontend_0i_115_13 (.A(frontend_0_n_115_8),.ZN(inst_src[4]));
	NAND2_X1_LVT frontend_0i_114_8 (.A1(frontend_0_n_114_6),.A2(frontend_0_n_114_7),.ZN(frontend_0_n_114_8));
	NOR2_X1_LVT frontend_0i_114_15 (.A1(frontend_0_n_114_5),.A2(frontend_0_n_114_8),.ZN(frontend_0_n_185));
	AOI22_X1_LVT frontend_0i_115_10 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_115),.B1(inst_type[2]),.B2(frontend_0_n_185),.ZN(frontend_0_n_115_7));
	INV_X1_LVT frontend_0i_115_11 (.A(frontend_0_n_115_7),.ZN(inst_src[3]));
	NOR2_X1_LVT frontend_0i_114_14 (.A1(frontend_0_n_114_4),.A2(frontend_0_n_114_8),.ZN(frontend_0_n_184));
	AOI22_X1_LVT frontend_0i_115_8 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_114),.B1(inst_type[2]),.B2(frontend_0_n_184),.ZN(frontend_0_n_115_6));
	INV_X1_LVT frontend_0i_115_9 (.A(frontend_0_n_115_6),.ZN(inst_src[2]));
	INV_X1_LVT frontend_0i_115_5 (.A(inst_type[2]),.ZN(frontend_0_n_115_4));
	NOR2_X1_LVT frontend_0i_114_13 (.A1(frontend_0_n_114_3),.A2(frontend_0_n_114_8),.ZN(frontend_0_n_183));
	AOI222_X1_LVT frontend_0i_115_6 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_113),.B1(frontend_0_n_115_4),.B2(inst_so[6]),.C1(inst_type[2]),.C2(frontend_0_n_183),.ZN(frontend_0_n_115_5));
	INV_X1_LVT frontend_0i_115_7 (.A(frontend_0_n_115_5),.ZN(inst_src[1]));
	NOR2_X1_LVT frontend_0i_114_12 (.A1(frontend_0_n_114_2),.A2(frontend_0_n_114_8),.ZN(frontend_0_n_182));
	AOI222_X1_LVT frontend_0i_115_3 (.A1(frontend_0_n_115_2),.A2(frontend_0_n_112),.B1(frontend_0_n_115_0),.B2(inst_so[7]),.C1(frontend_0_n_182),.C2(inst_type[2]),.ZN(frontend_0_n_115_3));
	INV_X1_LVT frontend_0i_115_4 (.A(frontend_0_n_115_3),.ZN(inst_src[0]));
	NOR3_X1_LVT frontend_0i_6_7 (.A1(frontend_0_i_state[0]),.A2(frontend_0_i_state[1]),.A3(frontend_0_i_state[2]),.ZN(frontend_0_n_8));
	NOR2_X1_LVT frontend_0i_118_0 (.A1(irq[13]),.A2(nmi_pnd),.ZN(frontend_0_n_118_0));
	INV_X1_LVT frontend_0i_118_1 (.A(frontend_0_n_118_0),.ZN(frontend_0_n_118_1));
	NOR2_X1_LVT frontend_0i_118_2 (.A1(frontend_0_n_118_1),.A2(irq[12]),.ZN(frontend_0_n_118_2));
	INV_X1_LVT frontend_0i_118_3 (.A(frontend_0_n_118_2),.ZN(frontend_0_n_118_3));
	NOR2_X1_LVT frontend_0i_118_4 (.A1(frontend_0_n_118_3),.A2(irq[11]),.ZN(frontend_0_n_118_4));
	INV_X1_LVT frontend_0i_118_5 (.A(frontend_0_n_118_4),.ZN(frontend_0_n_118_5));
	OR2_X1_LVT frontend_0i_116_0 (.A1(irq[10]),.A2(wdt_irq),.ZN(frontend_0_n_198));
	NOR2_X1_LVT frontend_0i_118_6 (.A1(frontend_0_n_118_5),.A2(frontend_0_n_198),.ZN(frontend_0_n_118_6));
	INV_X1_LVT frontend_0i_118_7 (.A(irq[9]),.ZN(frontend_0_n_118_7));
	NAND2_X1_LVT frontend_0i_118_8 (.A1(frontend_0_n_118_6),.A2(frontend_0_n_118_7),.ZN(frontend_0_n_118_8));
	NOR2_X1_LVT frontend_0i_118_9 (.A1(frontend_0_n_118_8),.A2(irq[8]),.ZN(frontend_0_n_118_9));
	INV_X1_LVT frontend_0i_118_10 (.A(frontend_0_n_118_9),.ZN(frontend_0_n_118_10));
	NOR2_X1_LVT frontend_0i_118_11 (.A1(frontend_0_n_118_10),.A2(irq[7]),.ZN(frontend_0_n_118_11));
	INV_X1_LVT frontend_0i_118_12 (.A(frontend_0_n_118_11),.ZN(frontend_0_n_118_12));
	NOR2_X1_LVT frontend_0i_118_13 (.A1(frontend_0_n_118_12),.A2(irq[6]),.ZN(frontend_0_n_118_13));
	INV_X1_LVT frontend_0i_118_14 (.A(irq[5]),.ZN(frontend_0_n_118_14));
	NAND2_X1_LVT frontend_0i_118_15 (.A1(frontend_0_n_118_13),.A2(frontend_0_n_118_14),.ZN(frontend_0_n_118_15));
	NOR2_X1_LVT frontend_0i_118_16 (.A1(frontend_0_n_118_15),.A2(irq[4]),.ZN(frontend_0_n_118_16));
	INV_X1_LVT frontend_0i_118_17 (.A(irq[3]),.ZN(frontend_0_n_118_17));
	NAND2_X1_LVT frontend_0i_118_18 (.A1(frontend_0_n_118_16),.A2(frontend_0_n_118_17),.ZN(frontend_0_n_118_18));
	NOR2_X1_LVT frontend_0i_118_19 (.A1(frontend_0_n_118_18),.A2(irq[2]),.ZN(frontend_0_n_118_19));
	NAND2_X1_LVT frontend_0i_118_20 (.A1(frontend_0_n_118_19),.A2(irq[1]),.ZN(frontend_0_n_118_20));
	INV_X1_LVT frontend_0i_118_21 (.A(frontend_0_n_118_20),.ZN(frontend_0_n_118_21));
	NAND2_X1_LVT frontend_0i_118_22 (.A1(frontend_0_n_118_9),.A2(irq[7]),.ZN(frontend_0_n_118_22));
	NAND2_X1_LVT frontend_0i_118_23 (.A1(frontend_0_n_118_6),.A2(irq[9]),.ZN(frontend_0_n_118_23));
	NAND2_X1_LVT frontend_0i_118_24 (.A1(frontend_0_n_118_2),.A2(irq[11]),.ZN(frontend_0_n_118_24));
	INV_X1_LVT frontend_0i_118_25 (.A(nmi_pnd),.ZN(frontend_0_n_118_25));
	NAND2_X1_LVT frontend_0i_118_26 (.A1(frontend_0_n_118_25),.A2(irq[13]),.ZN(frontend_0_n_118_26));
	NAND4_X1_LVT frontend_0i_118_27 (.A1(frontend_0_n_118_22),.A2(frontend_0_n_118_23),.A3(frontend_0_n_118_24),.A4(frontend_0_n_118_26),.ZN(frontend_0_n_118_27));
	AND2_X1_LVT frontend_0i_118_28 (.A1(frontend_0_n_118_16),.A2(irq[3]),.ZN(frontend_0_n_118_28));
	NAND2_X1_LVT frontend_0i_118_29 (.A1(frontend_0_n_118_13),.A2(irq[5]),.ZN(frontend_0_n_118_29));
	INV_X1_LVT frontend_0i_118_30 (.A(frontend_0_n_118_29),.ZN(frontend_0_n_118_30));
	NOR4_X1_LVT frontend_0i_118_31 (.A1(frontend_0_n_118_21),.A2(frontend_0_n_118_27),.A3(frontend_0_n_118_28),.A4(frontend_0_n_118_30),.ZN(frontend_0_n_118_31));
	INV_X1_LVT frontend_0i_118_32 (.A(frontend_0_n_118_19),.ZN(frontend_0_n_118_32));
	NOR2_X1_LVT frontend_0i_118_33 (.A1(frontend_0_n_118_32),.A2(irq[1]),.ZN(frontend_0_n_118_33));
	INV_X1_LVT frontend_0i_118_34 (.A(irq[0]),.ZN(frontend_0_n_118_34));
	NAND2_X1_LVT frontend_0i_118_35 (.A1(frontend_0_n_118_33),.A2(frontend_0_n_118_34),.ZN(frontend_0_n_118_35));
	NAND2_X1_LVT frontend_0i_118_36 (.A1(frontend_0_n_118_31),.A2(frontend_0_n_118_35),.ZN(frontend_0_n_200));
	CLKGATETST_X1_LVT frontend_0clk_gate_irq_num_reg (.CK(cpu_mclk),.E(frontend_0_irq_detect),.SE(1'b0),.GCK(frontend_0_n_199));
	DFFS_X1_LVT frontend_0irq_num_reg___05F05b0___05F05d (.D(frontend_0_n_200),.SN(frontend_0_n_91),.CK(frontend_0_n_199),.Q(frontend_0_irq_num[0]),.QN());
	INV_X1_LVT frontend_0i_120_0 (.A(frontend_0_irq_num[0]),.ZN(frontend_0_n_120_0));
	INV_X1_LVT frontend_0i_118_37 (.A(irq[2]),.ZN(frontend_0_n_118_36));
	NOR2_X1_LVT frontend_0i_118_38 (.A1(frontend_0_n_118_18),.A2(frontend_0_n_118_36),.ZN(frontend_0_n_118_37));
	NAND2_X1_LVT frontend_0i_118_39 (.A1(frontend_0_n_118_4),.A2(frontend_0_n_198),.ZN(frontend_0_n_118_38));
	NAND4_X1_LVT frontend_0i_118_40 (.A1(frontend_0_n_118_22),.A2(frontend_0_n_118_38),.A3(frontend_0_n_118_24),.A4(frontend_0_n_118_25),.ZN(frontend_0_n_118_39));
	NAND2_X1_LVT frontend_0i_118_41 (.A1(frontend_0_n_118_11),.A2(irq[6]),.ZN(frontend_0_n_118_40));
	INV_X1_LVT frontend_0i_118_42 (.A(frontend_0_n_118_40),.ZN(frontend_0_n_118_41));
	NOR4_X1_LVT frontend_0i_118_43 (.A1(frontend_0_n_118_37),.A2(frontend_0_n_118_39),.A3(frontend_0_n_118_28),.A4(frontend_0_n_118_41),.ZN(frontend_0_n_118_42));
	NAND2_X1_LVT frontend_0i_118_44 (.A1(frontend_0_n_118_42),.A2(frontend_0_n_118_35),.ZN(frontend_0_n_201));
	DFFS_X1_LVT frontend_0irq_num_reg___05F05b1___05F05d (.D(frontend_0_n_201),.SN(frontend_0_n_91),.CK(frontend_0_n_199),.Q(frontend_0_irq_num[1]),.QN());
	NOR2_X1_LVT frontend_0i_120_3 (.A1(frontend_0_n_120_0),.A2(frontend_0_irq_num[1]),.ZN(frontend_0_n_120_3));
	NAND2_X1_LVT frontend_0i_118_45 (.A1(frontend_0_n_118_0),.A2(irq[12]),.ZN(frontend_0_n_118_43));
	NAND4_X1_LVT frontend_0i_118_46 (.A1(frontend_0_n_118_22),.A2(frontend_0_n_118_43),.A3(frontend_0_n_118_26),.A4(frontend_0_n_118_25),.ZN(frontend_0_n_118_44));
	INV_X1_LVT frontend_0i_118_47 (.A(irq[4]),.ZN(frontend_0_n_118_45));
	NOR2_X1_LVT frontend_0i_118_48 (.A1(frontend_0_n_118_15),.A2(frontend_0_n_118_45),.ZN(frontend_0_n_118_46));
	NOR4_X1_LVT frontend_0i_118_49 (.A1(frontend_0_n_118_44),.A2(frontend_0_n_118_46),.A3(frontend_0_n_118_30),.A4(frontend_0_n_118_41),.ZN(frontend_0_n_118_47));
	NAND2_X1_LVT frontend_0i_118_50 (.A1(frontend_0_n_118_47),.A2(frontend_0_n_118_35),.ZN(frontend_0_n_202));
	DFFS_X1_LVT frontend_0irq_num_reg___05F05b2___05F05d (.D(frontend_0_n_202),.SN(frontend_0_n_91),.CK(frontend_0_n_199),.Q(frontend_0_irq_num[2]),.QN());
	NAND2_X1_LVT frontend_0i_120_12 (.A1(frontend_0_n_120_3),.A2(frontend_0_irq_num[2]),.ZN(frontend_0_n_120_12));
	NAND4_X1_LVT frontend_0i_118_51 (.A1(frontend_0_n_118_24),.A2(frontend_0_n_118_43),.A3(frontend_0_n_118_26),.A4(frontend_0_n_118_25),.ZN(frontend_0_n_118_48));
	INV_X1_LVT frontend_0i_118_52 (.A(irq[8]),.ZN(frontend_0_n_118_49));
	NOR2_X1_LVT frontend_0i_118_53 (.A1(frontend_0_n_118_8),.A2(frontend_0_n_118_49),.ZN(frontend_0_n_118_50));
	INV_X1_LVT frontend_0i_118_54 (.A(frontend_0_n_118_23),.ZN(frontend_0_n_118_51));
	INV_X1_LVT frontend_0i_118_55 (.A(frontend_0_n_118_38),.ZN(frontend_0_n_118_52));
	NOR4_X1_LVT frontend_0i_118_56 (.A1(frontend_0_n_118_48),.A2(frontend_0_n_118_50),.A3(frontend_0_n_118_51),.A4(frontend_0_n_118_52),.ZN(frontend_0_n_118_53));
	NAND2_X1_LVT frontend_0i_118_57 (.A1(frontend_0_n_118_53),.A2(frontend_0_n_118_35),.ZN(frontend_0_n_203));
	DFFS_X1_LVT frontend_0irq_num_reg___05F05b3___05F05d (.D(frontend_0_n_203),.SN(frontend_0_n_91),.CK(frontend_0_n_199),.Q(frontend_0_irq_num[3]),.QN());
	INV_X1_LVT frontend_0i_120_15 (.A(frontend_0_irq_num[3]),.ZN(frontend_0_n_120_15));
	NAND4_X1_LVT frontend_0i_118_58 (.A1(frontend_0_n_118_53),.A2(frontend_0_n_118_29),.A3(frontend_0_n_118_40),.A4(frontend_0_n_118_22),.ZN(frontend_0_n_118_54));
	NOR4_X1_LVT frontend_0i_118_59 (.A1(frontend_0_n_118_54),.A2(frontend_0_n_118_37),.A3(frontend_0_n_118_28),.A4(frontend_0_n_118_46),.ZN(frontend_0_n_118_55));
	NAND2_X1_LVT frontend_0i_118_60 (.A1(frontend_0_n_118_33),.A2(irq[0]),.ZN(frontend_0_n_118_56));
	NAND4_X1_LVT frontend_0i_118_61 (.A1(frontend_0_n_118_55),.A2(frontend_0_n_118_56),.A3(frontend_0_n_118_35),.A4(frontend_0_n_118_20),.ZN(frontend_0_n_204));
	DFFS_X1_LVT frontend_0irq_num_reg___05F05b4___05F05d (.D(frontend_0_n_204),.SN(frontend_0_n_91),.CK(frontend_0_n_199),.Q(frontend_0_irq_num[4]),.QN());
	INV_X1_LVT frontend_0i_120_16 (.A(frontend_0_irq_num[4]),.ZN(frontend_0_n_120_16));
	NOR2_X1_LVT frontend_0i_120_18 (.A1(frontend_0_n_120_15),.A2(frontend_0_n_120_16),.ZN(frontend_0_n_120_18));
	DFFS_X1_LVT frontend_0irq_num_reg___05F05b5___05F05d (.D(frontend_0_n_204),.SN(frontend_0_n_91),.CK(frontend_0_n_199),.Q(frontend_0_irq_num[5]),.QN());
	NAND2_X1_LVT frontend_0i_120_20 (.A1(frontend_0_n_120_18),.A2(frontend_0_irq_num[5]),.ZN(frontend_0_n_120_20));
	NOR2_X1_LVT frontend_0i_120_34 (.A1(frontend_0_n_120_12),.A2(frontend_0_n_120_20),.ZN(frontend_0_n_218));
	AND2_X1_LVT frontend_0i_121_13 (.A1(frontend_0_n_8),.A2(frontend_0_n_218),.ZN(irq_acc[13]));
	NOR2_X1_LVT frontend_0i_120_2 (.A1(frontend_0_irq_num[0]),.A2(frontend_0_irq_num[1]),.ZN(frontend_0_n_120_2));
	NAND2_X1_LVT frontend_0i_120_11 (.A1(frontend_0_n_120_2),.A2(frontend_0_irq_num[2]),.ZN(frontend_0_n_120_11));
	NOR2_X1_LVT frontend_0i_120_33 (.A1(frontend_0_n_120_11),.A2(frontend_0_n_120_20),.ZN(frontend_0_n_217));
	AND2_X1_LVT frontend_0i_121_12 (.A1(frontend_0_n_8),.A2(frontend_0_n_217),.ZN(irq_acc[12]));
	INV_X1_LVT frontend_0i_120_1 (.A(frontend_0_irq_num[1]),.ZN(frontend_0_n_120_1));
	NOR2_X1_LVT frontend_0i_120_5 (.A1(frontend_0_n_120_0),.A2(frontend_0_n_120_1),.ZN(frontend_0_n_120_5));
	INV_X1_LVT frontend_0i_120_6 (.A(frontend_0_irq_num[2]),.ZN(frontend_0_n_120_6));
	NAND2_X1_LVT frontend_0i_120_10 (.A1(frontend_0_n_120_5),.A2(frontend_0_n_120_6),.ZN(frontend_0_n_120_10));
	NOR2_X1_LVT frontend_0i_120_32 (.A1(frontend_0_n_120_10),.A2(frontend_0_n_120_20),.ZN(frontend_0_n_216));
	AND2_X1_LVT frontend_0i_121_11 (.A1(frontend_0_n_8),.A2(frontend_0_n_216),.ZN(irq_acc[11]));
	NOR2_X1_LVT frontend_0i_120_4 (.A1(frontend_0_irq_num[0]),.A2(frontend_0_n_120_1),.ZN(frontend_0_n_120_4));
	NAND2_X1_LVT frontend_0i_120_9 (.A1(frontend_0_n_120_4),.A2(frontend_0_n_120_6),.ZN(frontend_0_n_120_9));
	NOR2_X1_LVT frontend_0i_120_31 (.A1(frontend_0_n_120_9),.A2(frontend_0_n_120_20),.ZN(frontend_0_n_215));
	AND2_X1_LVT frontend_0i_121_10 (.A1(frontend_0_n_8),.A2(frontend_0_n_215),.ZN(irq_acc[10]));
	NAND2_X1_LVT frontend_0i_120_8 (.A1(frontend_0_n_120_3),.A2(frontend_0_n_120_6),.ZN(frontend_0_n_120_8));
	NOR2_X1_LVT frontend_0i_120_30 (.A1(frontend_0_n_120_8),.A2(frontend_0_n_120_20),.ZN(frontend_0_n_214));
	AND2_X1_LVT frontend_0i_121_9 (.A1(frontend_0_n_8),.A2(frontend_0_n_214),.ZN(irq_acc[9]));
	NAND2_X1_LVT frontend_0i_120_7 (.A1(frontend_0_n_120_2),.A2(frontend_0_n_120_6),.ZN(frontend_0_n_120_7));
	NOR2_X1_LVT frontend_0i_120_29 (.A1(frontend_0_n_120_7),.A2(frontend_0_n_120_20),.ZN(frontend_0_n_213));
	AND2_X1_LVT frontend_0i_121_8 (.A1(frontend_0_n_8),.A2(frontend_0_n_213),.ZN(irq_acc[8]));
	NAND2_X1_LVT frontend_0i_120_14 (.A1(frontend_0_n_120_5),.A2(frontend_0_irq_num[2]),.ZN(frontend_0_n_120_14));
	NOR2_X1_LVT frontend_0i_120_17 (.A1(frontend_0_irq_num[3]),.A2(frontend_0_n_120_16),.ZN(frontend_0_n_120_17));
	NAND2_X1_LVT frontend_0i_120_19 (.A1(frontend_0_n_120_17),.A2(frontend_0_irq_num[5]),.ZN(frontend_0_n_120_19));
	NOR2_X1_LVT frontend_0i_120_28 (.A1(frontend_0_n_120_14),.A2(frontend_0_n_120_19),.ZN(frontend_0_n_212));
	AND2_X1_LVT frontend_0i_121_7 (.A1(frontend_0_n_8),.A2(frontend_0_n_212),.ZN(irq_acc[7]));
	NAND2_X1_LVT frontend_0i_120_13 (.A1(frontend_0_n_120_4),.A2(frontend_0_irq_num[2]),.ZN(frontend_0_n_120_13));
	NOR2_X1_LVT frontend_0i_120_27 (.A1(frontend_0_n_120_13),.A2(frontend_0_n_120_19),.ZN(frontend_0_n_211));
	AND2_X1_LVT frontend_0i_121_6 (.A1(frontend_0_n_8),.A2(frontend_0_n_211),.ZN(irq_acc[6]));
	NOR2_X1_LVT frontend_0i_120_26 (.A1(frontend_0_n_120_12),.A2(frontend_0_n_120_19),.ZN(frontend_0_n_210));
	AND2_X1_LVT frontend_0i_121_5 (.A1(frontend_0_n_8),.A2(frontend_0_n_210),.ZN(irq_acc[5]));
	NOR2_X1_LVT frontend_0i_120_25 (.A1(frontend_0_n_120_11),.A2(frontend_0_n_120_19),.ZN(frontend_0_n_209));
	AND2_X1_LVT frontend_0i_121_4 (.A1(frontend_0_n_8),.A2(frontend_0_n_209),.ZN(irq_acc[4]));
	NOR2_X1_LVT frontend_0i_120_24 (.A1(frontend_0_n_120_10),.A2(frontend_0_n_120_19),.ZN(frontend_0_n_208));
	AND2_X1_LVT frontend_0i_121_3 (.A1(frontend_0_n_8),.A2(frontend_0_n_208),.ZN(irq_acc[3]));
	NOR2_X1_LVT frontend_0i_120_23 (.A1(frontend_0_n_120_9),.A2(frontend_0_n_120_19),.ZN(frontend_0_n_207));
	AND2_X1_LVT frontend_0i_121_2 (.A1(frontend_0_n_8),.A2(frontend_0_n_207),.ZN(irq_acc[2]));
	NOR2_X1_LVT frontend_0i_120_22 (.A1(frontend_0_n_120_8),.A2(frontend_0_n_120_19),.ZN(frontend_0_n_206));
	AND2_X1_LVT frontend_0i_121_1 (.A1(frontend_0_n_8),.A2(frontend_0_n_206),.ZN(irq_acc[1]));
	NOR2_X1_LVT frontend_0i_120_21 (.A1(frontend_0_n_120_7),.A2(frontend_0_n_120_19),.ZN(frontend_0_n_205));
	AND2_X1_LVT frontend_0i_121_0 (.A1(frontend_0_n_8),.A2(frontend_0_n_205),.ZN(irq_acc[0]));
	INV_X1_LVT frontend_0i_127_0 (.A(pc_sw_wr),.ZN(frontend_0_n_127_0));
	NOR3_X1_LVT frontend_0i_125_2 (.A1(frontend_0_i_state[0]),.A2(frontend_0_i_state[1]),.A3(frontend_0_i_state[2]),.ZN(frontend_0_n_221));
	INV_X1_LVT frontend_0i_125_0 (.A(frontend_0_i_state[0]),.ZN(frontend_0_n_125_0));
	NOR3_X1_LVT frontend_0i_125_1 (.A1(frontend_0_n_125_0),.A2(frontend_0_i_state[1]),.A3(frontend_0_i_state[2]),.ZN(frontend_0_n_220));
	NOR2_X1_LVT frontend_0i_125_3 (.A1(frontend_0_n_220),.A2(frontend_0_n_221),.ZN(frontend_0_n_222));
	DFFR_X1_LVT frontend_0pc_reg___05F05b15___05F05d (.D(pc_nxt[15]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[15]),.QN());
	AOI221_X1_LVT frontend_0i_126_28 (.A(frontend_0_n_221),.B1(frontend_0_n_220),.B2(fe_mdb_in[14]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[14]),.ZN(frontend_0_n_126_14));
	INV_X1_LVT frontend_0i_126_29 (.A(frontend_0_n_126_14),.ZN(frontend_0_n_237));
	AOI22_X1_LVT frontend_0i_127_29 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_237),.B1(pc_sw_wr),.B2(pc_sw[14]),.ZN(frontend_0_n_127_15));
	INV_X1_LVT frontend_0i_127_30 (.A(frontend_0_n_127_15),.ZN(pc_nxt[14]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b14___05F05d (.D(pc_nxt[14]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[14]),.QN());
	AOI221_X1_LVT frontend_0i_126_26 (.A(frontend_0_n_221),.B1(frontend_0_n_220),.B2(fe_mdb_in[13]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[13]),.ZN(frontend_0_n_126_13));
	INV_X1_LVT frontend_0i_126_27 (.A(frontend_0_n_126_13),.ZN(frontend_0_n_236));
	AOI22_X1_LVT frontend_0i_127_27 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_236),.B1(pc_sw_wr),.B2(pc_sw[13]),.ZN(frontend_0_n_127_14));
	INV_X1_LVT frontend_0i_127_28 (.A(frontend_0_n_127_14),.ZN(pc_nxt[13]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b13___05F05d (.D(pc_nxt[13]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[13]),.QN());
	AOI221_X1_LVT frontend_0i_126_24 (.A(frontend_0_n_221),.B1(frontend_0_n_220),.B2(fe_mdb_in[12]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[12]),.ZN(frontend_0_n_126_12));
	INV_X1_LVT frontend_0i_126_25 (.A(frontend_0_n_126_12),.ZN(frontend_0_n_235));
	AOI22_X1_LVT frontend_0i_127_25 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_235),.B1(pc_sw_wr),.B2(pc_sw[12]),.ZN(frontend_0_n_127_13));
	INV_X1_LVT frontend_0i_127_26 (.A(frontend_0_n_127_13),.ZN(pc_nxt[12]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b12___05F05d (.D(pc_nxt[12]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[12]),.QN());
	AOI221_X1_LVT frontend_0i_126_22 (.A(frontend_0_n_221),.B1(frontend_0_n_220),.B2(fe_mdb_in[11]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[11]),.ZN(frontend_0_n_126_11));
	INV_X1_LVT frontend_0i_126_23 (.A(frontend_0_n_126_11),.ZN(frontend_0_n_234));
	AOI22_X1_LVT frontend_0i_127_23 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_234),.B1(pc_sw_wr),.B2(pc_sw[11]),.ZN(frontend_0_n_127_12));
	INV_X1_LVT frontend_0i_127_24 (.A(frontend_0_n_127_12),.ZN(pc_nxt[11]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b11___05F05d (.D(pc_nxt[11]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[11]),.QN());
	AOI221_X1_LVT frontend_0i_126_20 (.A(frontend_0_n_221),.B1(frontend_0_n_220),.B2(fe_mdb_in[10]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[10]),.ZN(frontend_0_n_126_10));
	INV_X1_LVT frontend_0i_126_21 (.A(frontend_0_n_126_10),.ZN(frontend_0_n_233));
	AOI22_X1_LVT frontend_0i_127_21 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_233),.B1(pc_sw_wr),.B2(pc_sw[10]),.ZN(frontend_0_n_127_11));
	INV_X1_LVT frontend_0i_127_22 (.A(frontend_0_n_127_11),.ZN(pc_nxt[10]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b10___05F05d (.D(pc_nxt[10]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[10]),.QN());
	AOI221_X1_LVT frontend_0i_126_18 (.A(frontend_0_n_221),.B1(frontend_0_n_220),.B2(fe_mdb_in[9]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[9]),.ZN(frontend_0_n_126_9));
	INV_X1_LVT frontend_0i_126_19 (.A(frontend_0_n_126_9),.ZN(frontend_0_n_232));
	AOI22_X1_LVT frontend_0i_127_19 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_232),.B1(pc_sw_wr),.B2(pc_sw[9]),.ZN(frontend_0_n_127_10));
	INV_X1_LVT frontend_0i_127_20 (.A(frontend_0_n_127_10),.ZN(pc_nxt[9]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b9___05F05d (.D(pc_nxt[9]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[9]),.QN());
	AOI221_X1_LVT frontend_0i_126_16 (.A(frontend_0_n_221),.B1(frontend_0_n_220),.B2(fe_mdb_in[8]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[8]),.ZN(frontend_0_n_126_8));
	INV_X1_LVT frontend_0i_126_17 (.A(frontend_0_n_126_8),.ZN(frontend_0_n_231));
	AOI22_X1_LVT frontend_0i_127_17 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_231),.B1(pc_sw_wr),.B2(pc_sw[8]),.ZN(frontend_0_n_127_9));
	INV_X1_LVT frontend_0i_127_18 (.A(frontend_0_n_127_9),.ZN(pc_nxt[8]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b8___05F05d (.D(pc_nxt[8]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[8]),.QN());
	AOI221_X1_LVT frontend_0i_126_14 (.A(frontend_0_n_221),.B1(frontend_0_n_220),.B2(fe_mdb_in[7]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[7]),.ZN(frontend_0_n_126_7));
	INV_X1_LVT frontend_0i_126_15 (.A(frontend_0_n_126_7),.ZN(frontend_0_n_230));
	AOI22_X1_LVT frontend_0i_127_15 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_230),.B1(pc_sw_wr),.B2(pc_sw[7]),.ZN(frontend_0_n_127_8));
	INV_X1_LVT frontend_0i_127_16 (.A(frontend_0_n_127_8),.ZN(pc_nxt[7]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b7___05F05d (.D(pc_nxt[7]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[7]),.QN());
	AOI222_X1_LVT frontend_0i_126_12 (.A1(frontend_0_n_221),.A2(frontend_0_irq_num[5]),.B1(frontend_0_n_220),.B2(fe_mdb_in[6]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[6]),.ZN(frontend_0_n_126_6));
	INV_X1_LVT frontend_0i_126_13 (.A(frontend_0_n_126_6),.ZN(frontend_0_n_229));
	AOI22_X1_LVT frontend_0i_127_13 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_229),.B1(pc_sw_wr),.B2(pc_sw[6]),.ZN(frontend_0_n_127_7));
	INV_X1_LVT frontend_0i_127_14 (.A(frontend_0_n_127_7),.ZN(pc_nxt[6]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b6___05F05d (.D(pc_nxt[6]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[6]),.QN());
	AOI222_X1_LVT frontend_0i_126_10 (.A1(frontend_0_n_221),.A2(frontend_0_irq_num[4]),.B1(frontend_0_n_220),.B2(fe_mdb_in[5]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[5]),.ZN(frontend_0_n_126_5));
	INV_X1_LVT frontend_0i_126_11 (.A(frontend_0_n_126_5),.ZN(frontend_0_n_228));
	AOI22_X1_LVT frontend_0i_127_11 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_228),.B1(pc_sw_wr),.B2(pc_sw[5]),.ZN(frontend_0_n_127_6));
	INV_X1_LVT frontend_0i_127_12 (.A(frontend_0_n_127_6),.ZN(pc_nxt[5]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b5___05F05d (.D(pc_nxt[5]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[5]),.QN());
	AOI222_X1_LVT frontend_0i_126_8 (.A1(frontend_0_n_221),.A2(frontend_0_irq_num[3]),.B1(frontend_0_n_220),.B2(fe_mdb_in[4]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[4]),.ZN(frontend_0_n_126_4));
	INV_X1_LVT frontend_0i_126_9 (.A(frontend_0_n_126_4),.ZN(frontend_0_n_227));
	AOI22_X1_LVT frontend_0i_127_9 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_227),.B1(pc_sw_wr),.B2(pc_sw[4]),.ZN(frontend_0_n_127_5));
	INV_X1_LVT frontend_0i_127_10 (.A(frontend_0_n_127_5),.ZN(pc_nxt[4]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b4___05F05d (.D(pc_nxt[4]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[4]),.QN());
	AOI222_X1_LVT frontend_0i_126_6 (.A1(frontend_0_n_221),.A2(frontend_0_irq_num[2]),.B1(frontend_0_n_220),.B2(fe_mdb_in[3]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[3]),.ZN(frontend_0_n_126_3));
	INV_X1_LVT frontend_0i_126_7 (.A(frontend_0_n_126_3),.ZN(frontend_0_n_226));
	AOI22_X1_LVT frontend_0i_127_7 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_226),.B1(pc_sw_wr),.B2(pc_sw[3]),.ZN(frontend_0_n_127_4));
	INV_X1_LVT frontend_0i_127_8 (.A(frontend_0_n_127_4),.ZN(pc_nxt[3]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b3___05F05d (.D(pc_nxt[3]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[3]),.QN());
	AOI222_X1_LVT frontend_0i_126_4 (.A1(frontend_0_n_221),.A2(frontend_0_irq_num[1]),.B1(frontend_0_n_220),.B2(fe_mdb_in[2]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[2]),.ZN(frontend_0_n_126_2));
	INV_X1_LVT frontend_0i_126_5 (.A(frontend_0_n_126_2),.ZN(frontend_0_n_225));
	AOI22_X1_LVT frontend_0i_127_5 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_225),.B1(pc_sw_wr),.B2(pc_sw[2]),.ZN(frontend_0_n_127_3));
	INV_X1_LVT frontend_0i_127_6 (.A(frontend_0_n_127_3),.ZN(pc_nxt[2]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b2___05F05d (.D(pc_nxt[2]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[2]),.QN());
	INV_X1_LVT frontend_0i_122_0 (.A(frontend_0_e_state_nxt_reg[1]),.ZN(frontend_0_n_122_0));
	AND4_X1_LVT frontend_0i_122_1 (.A1(frontend_0_n_122_0),.A2(frontend_0_e_state_nxt_reg[0]),.A3(frontend_0_e_state_nxt_reg[2]),.A4(frontend_0_e_state_nxt_reg[3]),.ZN(frontend_0_n_122_1));
	INV_X1_LVT frontend_0i_122_2 (.A(frontend_0_n_73),.ZN(frontend_0_n_122_2));
	AOI21_X1_LVT frontend_0i_122_3 (.A(frontend_0_n_122_1),.B1(frontend_0_n_122_2),.B2(frontend_0_n_4),.ZN(frontend_0_fetch));
	AOI222_X1_LVT frontend_0i_126_2 (.A1(frontend_0_n_221),.A2(frontend_0_irq_num[0]),.B1(frontend_0_n_220),.B2(fe_mdb_in[1]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[1]),.ZN(frontend_0_n_126_1));
	INV_X1_LVT frontend_0i_126_3 (.A(frontend_0_n_126_1),.ZN(frontend_0_n_224));
	AOI22_X1_LVT frontend_0i_127_3 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_224),.B1(pc_sw_wr),.B2(pc_sw[1]),.ZN(frontend_0_n_127_2));
	INV_X1_LVT frontend_0i_127_4 (.A(frontend_0_n_127_2),.ZN(pc_nxt[1]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b1___05F05d (.D(pc_nxt[1]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[1]),.QN());
	HA_X1_LVT frontend_0i_124_0 (.A(frontend_0_fetch),.B(pc[1]),.CO(frontend_0_n_124_0),.S(frontend_0_pc_incr[1]));
	HA_X1_LVT frontend_0i_124_1 (.A(pc[2]),.B(frontend_0_n_124_0),.CO(frontend_0_n_124_1),.S(frontend_0_pc_incr[2]));
	HA_X1_LVT frontend_0i_124_2 (.A(pc[3]),.B(frontend_0_n_124_1),.CO(frontend_0_n_124_2),.S(frontend_0_pc_incr[3]));
	HA_X1_LVT frontend_0i_124_3 (.A(pc[4]),.B(frontend_0_n_124_2),.CO(frontend_0_n_124_3),.S(frontend_0_pc_incr[4]));
	HA_X1_LVT frontend_0i_124_4 (.A(pc[5]),.B(frontend_0_n_124_3),.CO(frontend_0_n_124_4),.S(frontend_0_pc_incr[5]));
	HA_X1_LVT frontend_0i_124_5 (.A(pc[6]),.B(frontend_0_n_124_4),.CO(frontend_0_n_124_5),.S(frontend_0_pc_incr[6]));
	HA_X1_LVT frontend_0i_124_6 (.A(pc[7]),.B(frontend_0_n_124_5),.CO(frontend_0_n_124_6),.S(frontend_0_pc_incr[7]));
	HA_X1_LVT frontend_0i_124_7 (.A(pc[8]),.B(frontend_0_n_124_6),.CO(frontend_0_n_124_7),.S(frontend_0_pc_incr[8]));
	HA_X1_LVT frontend_0i_124_8 (.A(pc[9]),.B(frontend_0_n_124_7),.CO(frontend_0_n_124_8),.S(frontend_0_pc_incr[9]));
	HA_X1_LVT frontend_0i_124_9 (.A(pc[10]),.B(frontend_0_n_124_8),.CO(frontend_0_n_124_9),.S(frontend_0_pc_incr[10]));
	HA_X1_LVT frontend_0i_124_10 (.A(pc[11]),.B(frontend_0_n_124_9),.CO(frontend_0_n_124_10),.S(frontend_0_pc_incr[11]));
	HA_X1_LVT frontend_0i_124_11 (.A(pc[12]),.B(frontend_0_n_124_10),.CO(frontend_0_n_124_11),.S(frontend_0_pc_incr[12]));
	HA_X1_LVT frontend_0i_124_12 (.A(pc[13]),.B(frontend_0_n_124_11),.CO(frontend_0_n_124_12),.S(frontend_0_pc_incr[13]));
	HA_X1_LVT frontend_0i_124_13 (.A(pc[14]),.B(frontend_0_n_124_12),.CO(frontend_0_n_124_13),.S(frontend_0_pc_incr[14]));
	XNOR2_X1_LVT frontend_0i_124_14 (.A(pc[15]),.B(frontend_0_n_124_13),.ZN(frontend_0_n_124_14));
	INV_X1_LVT frontend_0i_124_15 (.A(frontend_0_n_124_14),.ZN(frontend_0_pc_incr[15]));
	AOI221_X1_LVT frontend_0i_126_30 (.A(frontend_0_n_221),.B1(frontend_0_n_220),.B2(fe_mdb_in[15]),.C1(frontend_0_n_222),.C2(frontend_0_pc_incr[15]),.ZN(frontend_0_n_126_15));
	INV_X1_LVT frontend_0i_126_31 (.A(frontend_0_n_126_15),.ZN(frontend_0_n_238));
	AOI22_X1_LVT frontend_0i_127_31 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_238),.B1(pc_sw_wr),.B2(pc_sw[15]),.ZN(frontend_0_n_127_16));
	INV_X1_LVT frontend_0i_127_32 (.A(frontend_0_n_127_16),.ZN(pc_nxt[15]));
	DFFR_X1_LVT frontend_0pc_reg___05F05b0___05F05d (.D(pc_nxt[0]),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(pc[0]),.QN());
	AOI22_X1_LVT frontend_0i_126_0 (.A1(fe_mdb_in[0]),.A2(frontend_0_n_220),.B1(pc[0]),.B2(frontend_0_n_222),.ZN(frontend_0_n_126_0));
	INV_X1_LVT frontend_0i_126_1 (.A(frontend_0_n_126_0),.ZN(frontend_0_n_223));
	AOI22_X1_LVT frontend_0i_127_1 (.A1(frontend_0_n_127_0),.A2(frontend_0_n_223),.B1(pc_sw[0]),.B2(pc_sw_wr),.ZN(frontend_0_n_127_1));
	INV_X1_LVT frontend_0i_127_2 (.A(frontend_0_n_127_1),.ZN(pc_nxt[0]));
	DFFR_X1_LVT frontend_0pmem_busy_reg (.D(fe_pmem_wait),.RN(frontend_0_n_91),.CK(cpu_mclk),.Q(frontend_0_pmem_busy),.QN());
	NOR4_X1_LVT frontend_0i_128_0 (.A1(pc_sw_wr),.A2(frontend_0_fetch),.A3(frontend_0_pmem_busy),.A4(frontend_0_n_8),.ZN(frontend_0_n_128_0));
	NAND2_X1_LVT frontend_0i_128_1 (.A1(cpu_halt_st),.A2(frontend_0_n_0),.ZN(frontend_0_n_128_1));
	NAND2_X1_LVT frontend_0i_128_2 (.A1(frontend_0_n_128_0),.A2(frontend_0_n_128_1),.ZN(fe_mb_en));
	AND2_X1_LVT frontend_0i_129_0 (.A1(dma_en),.A2(cpu_en_s),.ZN(mclk_dma_enable));
	AND2_X1_LVT frontend_0and_mclk_dma_wkupi_0_0 (.A1(dma_wkup),.A2(cpu_en_s),.ZN(mclk_dma_wkup));
	INV_X1_LVT frontend_0i_130_0 (.A(cpu_en_s),.ZN(frontend_0_n_130_0));
	OAI211_X1_LVT frontend_0i_130_1 (.A(frontend_0_n_5),.B(frontend_0_n_67),.C1(frontend_0_n_130_0),.C2(cpuoff),.ZN(frontend_0_n_130_1));
	INV_X1_LVT frontend_0i_130_2 (.A(inst_irq_rst),.ZN(frontend_0_n_130_2));
	AOI22_X1_LVT frontend_0i_130_3 (.A1(frontend_0_n_130_1),.A2(frontend_0_n_130_2),.B1(cpu_en_s),.B2(inst_irq_rst),.ZN(frontend_0_n_130_3));
	INV_X1_LVT frontend_0i_130_4 (.A(frontend_0_n_130_3),.ZN(mclk_enable));
	OR2_X1_LVT frontend_0i_132_0 (.A1(wkup),.A2(wdt_wkup),.ZN(frontend_0_n_240));
	AND2_X1_LVT frontend_0and_mirq_wkupi_0_0 (.A1(frontend_0_n_240),.A2(gie),.ZN(frontend_0_mirq_wkup));
	OR2_X1_LVT frontend_0i_131_0 (.A1(nmi_wkup),.A2(frontend_0_mirq_wkup),.ZN(frontend_0_n_239));
	AND2_X1_LVT frontend_0and_mclk_wkupi_0_0 (.A1(frontend_0_n_239),.A2(cpu_en_s),.ZN(mclk_wkup));
	NOR2_X1_LVT frontend_0i_120_35 (.A1(frontend_0_n_120_13),.A2(frontend_0_n_120_20),.ZN(frontend_0_n_219));
	AND2_X1_LVT frontend_0i_121_14 (.A1(frontend_0_n_8),.A2(frontend_0_n_219),.ZN(nmi_acc));
	INV_X1_LVT execution_unit_0i_0_0 (.A(e_state[3]),.ZN(execution_unit_0_n_0_0));
	INV_X1_LVT execution_unit_0i_0_1 (.A(e_state[0]),.ZN(execution_unit_0_n_0_1));
	INV_X1_LVT execution_unit_0i_0_2 (.A(e_state[1]),.ZN(execution_unit_0_n_0_2));
	NOR4_X1_LVT execution_unit_0i_0_3 (.A1(execution_unit_0_n_0_0),.A2(execution_unit_0_n_0_1),.A3(execution_unit_0_n_0_2),.A4(e_state[2]),.ZN(execution_unit_0_n_0));
	OR3_X1_LVT execution_unit_0i_38_0 (.A1(inst_as[4]),.A2(inst_as[1]),.A3(inst_as[6]),.ZN(execution_unit_0_n_69));
	INV_X1_LVT execution_unit_0i_0_4 (.A(e_state[2]),.ZN(execution_unit_0_n_0_3));
	NOR4_X1_LVT execution_unit_0i_0_5 (.A1(execution_unit_0_n_0_2),.A2(execution_unit_0_n_0_3),.A3(e_state[0]),.A4(e_state[3]),.ZN(execution_unit_0_n_1));
	NOR4_X1_LVT execution_unit_0i_0_6 (.A1(execution_unit_0_n_0_3),.A2(execution_unit_0_n_0_1),.A3(execution_unit_0_n_0_2),.A4(e_state[3]),.ZN(execution_unit_0_n_2));
	AOI22_X1_LVT execution_unit_0i_39_11 (.A1(execution_unit_0_n_69),.A2(execution_unit_0_n_1),.B1(execution_unit_0_n_69),.B2(execution_unit_0_n_2),.ZN(execution_unit_0_n_39_8));
	INV_X1_LVT execution_unit_0i_39_12 (.A(execution_unit_0_n_39_8),.ZN(execution_unit_0_n_73));
	INV_X1_LVT execution_unit_0i_40_4 (.A(execution_unit_0_n_73),.ZN(execution_unit_0_n_40_4));
	NOR2_X1_LVT execution_unit_0i_40_5 (.A1(execution_unit_0_n_40_4),.A2(cpu_halt_st),.ZN(execution_unit_0_n_74));
	NAND2_X1_LVT execution_unit_0i_41_90 (.A1(execution_unit_0_n_74),.A2(inst_sext[15]),.ZN(execution_unit_0_n_41_75));
	OR2_X1_LVT execution_unit_0i_40_0 (.A1(execution_unit_0_n_73),.A2(cpu_halt_st),.ZN(execution_unit_0_n_40_0));
	NOR4_X1_LVT execution_unit_0i_0_7 (.A1(execution_unit_0_n_0_2),.A2(execution_unit_0_n_0_0),.A3(e_state[0]),.A4(e_state[2]),.ZN(execution_unit_0_n_3));
	AND2_X1_LVT execution_unit_0i_22_0 (.A1(inst_so[6]),.A2(execution_unit_0_n_3),.ZN(execution_unit_0_n_40));
	INV_X1_LVT execution_unit_0i_39_8 (.A(execution_unit_0_n_40),.ZN(execution_unit_0_n_39_6));
	INV_X1_LVT execution_unit_0i_2_0 (.A(inst_so[6]),.ZN(execution_unit_0_n_10));
	AND2_X1_LVT execution_unit_0i_36_0 (.A1(execution_unit_0_n_0),.A2(execution_unit_0_n_10),.ZN(execution_unit_0_n_67));
	INV_X1_LVT execution_unit_0i_39_9 (.A(execution_unit_0_n_67),.ZN(execution_unit_0_n_39_7));
	OR3_X1_LVT execution_unit_0i_37_0 (.A1(inst_ad[0]),.A2(inst_type[0]),.A3(inst_type[1]),.ZN(execution_unit_0_n_68));
	OAI21_X1_LVT execution_unit_0i_39_10 (.A(execution_unit_0_n_39_6),.B1(execution_unit_0_n_39_7),.B2(execution_unit_0_n_68),.ZN(execution_unit_0_n_72));
	INV_X1_LVT execution_unit_0i_40_6 (.A(execution_unit_0_n_72),.ZN(execution_unit_0_n_40_5));
	NOR2_X1_LVT execution_unit_0i_40_7 (.A1(execution_unit_0_n_40_0),.A2(execution_unit_0_n_40_5),.ZN(execution_unit_0_n_75));
	INV_X1_LVT execution_unit_0i_33_0 (.A(inst_bw),.ZN(execution_unit_0_n_47));
	INV_X1_LVT execution_unit_0i_6_0 (.A(inst_alu[11]),.ZN(execution_unit_0_n_13));
	INV_X1_LVT execution_unit_0i_3_0 (.A(inst_irq_rst),.ZN(execution_unit_0_n_11));
	NOR4_X1_LVT execution_unit_0i_0_10 (.A1(execution_unit_0_n_0_1),.A2(execution_unit_0_n_0_2),.A3(e_state[2]),.A4(e_state[3]),.ZN(execution_unit_0_n_6));
	NOR4_X1_LVT execution_unit_0i_0_9 (.A1(execution_unit_0_n_0_1),.A2(e_state[1]),.A3(e_state[2]),.A4(e_state[3]),.ZN(execution_unit_0_n_5));
	OAI21_X1_LVT execution_unit_0i_4_0 (.A(execution_unit_0_n_11),.B1(execution_unit_0_n_6),.B2(execution_unit_0_n_5),.ZN(execution_unit_0_n_4_0));
	NAND2_X1_LVT execution_unit_0i_4_1 (.A1(execution_unit_0_n_10),.A2(execution_unit_0_n_3),.ZN(execution_unit_0_n_4_1));
	NAND2_X1_LVT execution_unit_0i_4_2 (.A1(execution_unit_0_n_4_0),.A2(execution_unit_0_n_4_1),.ZN(execution_unit_0_n_12));
	OR2_X1_LVT execution_unit_0i_5_0 (.A1(execution_unit_0_n_12),.A2(execution_unit_0_n_2),.ZN(execution_unit_0_mb_wr_det));
	AND2_X1_LVT execution_unit_0i_7_0 (.A1(execution_unit_0_n_13),.A2(execution_unit_0_mb_wr_det),.ZN(execution_unit_0_n_7_0));
	NOR4_X1_LVT execution_unit_0i_0_8 (.A1(execution_unit_0_n_0_1),.A2(execution_unit_0_n_0_0),.A3(e_state[1]),.A4(e_state[2]),.ZN(execution_unit_0_n_4));
	INV_X1_LVT execution_unit_0i_7_1 (.A(execution_unit_0_n_4),.ZN(execution_unit_0_n_7_1));
	NOR3_X1_LVT execution_unit_0i_7_2 (.A1(execution_unit_0_n_7_1),.A2(inst_type[0]),.A3(inst_mov),.ZN(execution_unit_0_n_7_2));
	INV_X1_LVT execution_unit_0i_7_3 (.A(execution_unit_0_n_1),.ZN(execution_unit_0_n_7_3));
	NOR2_X1_LVT execution_unit_0i_7_4 (.A1(execution_unit_0_n_7_3),.A2(inst_as[5]),.ZN(execution_unit_0_n_7_4));
	AND2_X1_LVT execution_unit_0i_1_0 (.A1(execution_unit_0_n_0),.A2(inst_so[6]),.ZN(execution_unit_0_n_9));
	OR4_X1_LVT execution_unit_0i_7_5 (.A1(execution_unit_0_n_7_0),.A2(execution_unit_0_n_7_2),.A3(execution_unit_0_n_7_4),.A4(execution_unit_0_n_9),.ZN(eu_mb_en));
	CLKGATETST_X1_LVT execution_unit_0clk_gate_mab_lsb_reg (.CK(cpu_mclk),.E(eu_mb_en),.SE(1'b0),.GCK(execution_unit_0_n_16));
	INV_X1_LVT execution_unit_0i_11_0 (.A(puc_rst),.ZN(execution_unit_0_n_18));
	DFFR_X1_LVT execution_unit_0mab_lsb_reg (.D(eu_mab[0]),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_16),.Q(execution_unit_0_mab_lsb),.QN());
	AND2_X1_LVT execution_unit_0i_33_2 (.A1(execution_unit_0_mab_lsb),.A2(inst_bw),.ZN(execution_unit_0_n_49));
	NOR2_X1_LVT execution_unit_0i_33_1 (.A1(execution_unit_0_n_47),.A2(execution_unit_0_mab_lsb),.ZN(execution_unit_0_n_48));
	NOR3_X1_LVT execution_unit_0i_34_17 (.A1(execution_unit_0_n_47),.A2(execution_unit_0_n_49),.A3(execution_unit_0_n_48),.ZN(execution_unit_0_n_34_9));
	INV_X1_LVT execution_unit_0i_34_32 (.A(eu_mdb_in[15]),.ZN(execution_unit_0_n_34_17));
	NOR2_X1_LVT execution_unit_0i_34_33 (.A1(execution_unit_0_n_34_9),.A2(execution_unit_0_n_34_17),.ZN(execution_unit_0_n_65));
	NAND2_X1_LVT execution_unit_0i_41_91 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_65),.ZN(execution_unit_0_n_41_76));
	NOR2_X1_LVT execution_unit_0i_40_1 (.A1(execution_unit_0_n_40_0),.A2(execution_unit_0_n_72),.ZN(execution_unit_0_n_40_1));
	INV_X1_LVT execution_unit_0i_39_3 (.A(execution_unit_0_n_4),.ZN(execution_unit_0_n_39_2));
	OR2_X1_LVT execution_unit_0i_18_0 (.A1(inst_so[4]),.A2(inst_so[5]),.ZN(execution_unit_0_n_37));
	OR2_X1_LVT execution_unit_0i_19_0 (.A1(inst_so[6]),.A2(execution_unit_0_n_37),.ZN(execution_unit_0_n_38));
	NOR3_X1_LVT execution_unit_0i_39_4 (.A1(execution_unit_0_n_39_2),.A2(inst_ad[6]),.A3(execution_unit_0_n_38),.ZN(execution_unit_0_n_39_3));
	INV_X1_LVT execution_unit_0i_39_5 (.A(inst_ad[6]),.ZN(execution_unit_0_n_39_4));
	AOI221_X1_LVT execution_unit_0i_39_6 (.A(execution_unit_0_n_39_3),.B1(execution_unit_0_n_39_4),.B2(execution_unit_0_n_3),.C1(execution_unit_0_n_68),.C2(execution_unit_0_n_67),.ZN(execution_unit_0_n_39_5));
	INV_X1_LVT execution_unit_0i_39_7 (.A(execution_unit_0_n_39_5),.ZN(execution_unit_0_n_71));
	AND2_X1_LVT execution_unit_0i_40_8 (.A1(execution_unit_0_n_40_1),.A2(execution_unit_0_n_71),.ZN(execution_unit_0_n_76));
	NAND2_X1_LVT execution_unit_0i_41_92 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[15]),.ZN(execution_unit_0_n_41_77));
	INV_X1_LVT execution_unit_0i_40_2 (.A(execution_unit_0_n_71),.ZN(execution_unit_0_n_40_2));
	NAND2_X1_LVT execution_unit_0i_40_3 (.A1(execution_unit_0_n_40_1),.A2(execution_unit_0_n_40_2),.ZN(execution_unit_0_n_40_3));
	OR2_X1_LVT execution_unit_0i_24_0 (.A1(inst_as[2]),.A2(inst_as[3]),.ZN(execution_unit_0_n_41));
	AND2_X1_LVT execution_unit_0i_25_0 (.A1(inst_src[1]),.A2(execution_unit_0_n_41),.ZN(execution_unit_0_n_42));
	AND3_X1_LVT execution_unit_0i_26_0 (.A1(execution_unit_0_n_42),.A2(execution_unit_0_n_1),.A3(execution_unit_0_n_37),.ZN(execution_unit_0_n_43));
	NOR4_X1_LVT execution_unit_0i_0_12 (.A1(execution_unit_0_n_0_1),.A2(execution_unit_0_n_0_3),.A3(e_state[1]),.A4(e_state[3]),.ZN(execution_unit_0_n_8));
	AND3_X1_LVT execution_unit_0i_27_0 (.A1(inst_as[1]),.A2(execution_unit_0_n_8),.A3(execution_unit_0_n_37),.ZN(execution_unit_0_n_44));
	OR2_X1_LVT execution_unit_0i_29_0 (.A1(execution_unit_0_n_5),.A2(execution_unit_0_n_6),.ZN(execution_unit_0_n_46));
	OR2_X1_LVT execution_unit_0i_35_0 (.A1(execution_unit_0_n_44),.A2(execution_unit_0_n_46),.ZN(execution_unit_0_n_66));
	NOR4_X1_LVT execution_unit_0i_0_11 (.A1(execution_unit_0_n_0_2),.A2(e_state[0]),.A3(e_state[2]),.A4(e_state[3]),.ZN(execution_unit_0_n_7));
	NOR3_X1_LVT execution_unit_0i_39_0 (.A1(execution_unit_0_n_43),.A2(execution_unit_0_n_66),.A3(execution_unit_0_n_7),.ZN(execution_unit_0_n_39_0));
	AND2_X1_LVT execution_unit_0i_28_0 (.A1(execution_unit_0_n_37),.A2(execution_unit_0_n_4),.ZN(execution_unit_0_n_45));
	NAND2_X1_LVT execution_unit_0i_39_1 (.A1(execution_unit_0_n_10),.A2(execution_unit_0_n_45),.ZN(execution_unit_0_n_39_1));
	NAND2_X1_LVT execution_unit_0i_39_2 (.A1(execution_unit_0_n_39_0),.A2(execution_unit_0_n_39_1),.ZN(execution_unit_0_n_70));
	INV_X1_LVT execution_unit_0i_40_9 (.A(execution_unit_0_n_70),.ZN(execution_unit_0_n_40_6));
	NOR2_X1_LVT execution_unit_0i_40_10 (.A1(execution_unit_0_n_40_3),.A2(execution_unit_0_n_40_6),.ZN(execution_unit_0_n_77));
	INV_X1_LVT execution_unit_0i_41_8 (.A(execution_unit_0_n_77),.ZN(execution_unit_0_n_41_7));
	NAND4_X1_LVT execution_unit_0i_41_93 (.A1(execution_unit_0_n_41_75),.A2(execution_unit_0_n_41_76),.A3(execution_unit_0_n_41_77),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_78));
	AOI21_X1_LVT execution_unit_0i_41_94 (.A(execution_unit_0_n_41_78),.B1(cpu_halt_st),.B2(dbg_mem_dout[15]),.ZN(execution_unit_0_n_41_79));
	INV_X1_LVT execution_unit_0i_41_95 (.A(execution_unit_0_n_41_79),.ZN(execution_unit_0_n_93));
	NAND2_X1_LVT execution_unit_0i_41_84 (.A1(execution_unit_0_n_74),.A2(inst_sext[14]),.ZN(execution_unit_0_n_41_70));
	INV_X1_LVT execution_unit_0i_34_30 (.A(eu_mdb_in[14]),.ZN(execution_unit_0_n_34_16));
	NOR2_X1_LVT execution_unit_0i_34_31 (.A1(execution_unit_0_n_34_9),.A2(execution_unit_0_n_34_16),.ZN(execution_unit_0_n_64));
	NAND2_X1_LVT execution_unit_0i_41_85 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_64),.ZN(execution_unit_0_n_41_71));
	NAND2_X1_LVT execution_unit_0i_41_86 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[14]),.ZN(execution_unit_0_n_41_72));
	NAND4_X1_LVT execution_unit_0i_41_87 (.A1(execution_unit_0_n_41_70),.A2(execution_unit_0_n_41_71),.A3(execution_unit_0_n_41_72),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_73));
	AOI21_X1_LVT execution_unit_0i_41_88 (.A(execution_unit_0_n_41_73),.B1(cpu_halt_st),.B2(dbg_mem_dout[14]),.ZN(execution_unit_0_n_41_74));
	INV_X1_LVT execution_unit_0i_41_89 (.A(execution_unit_0_n_41_74),.ZN(execution_unit_0_n_92));
	NAND2_X1_LVT execution_unit_0i_41_78 (.A1(execution_unit_0_n_74),.A2(inst_sext[13]),.ZN(execution_unit_0_n_41_65));
	INV_X1_LVT execution_unit_0i_34_28 (.A(eu_mdb_in[13]),.ZN(execution_unit_0_n_34_15));
	NOR2_X1_LVT execution_unit_0i_34_29 (.A1(execution_unit_0_n_34_9),.A2(execution_unit_0_n_34_15),.ZN(execution_unit_0_n_63));
	NAND2_X1_LVT execution_unit_0i_41_79 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_63),.ZN(execution_unit_0_n_41_66));
	NAND2_X1_LVT execution_unit_0i_41_80 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[13]),.ZN(execution_unit_0_n_41_67));
	NAND4_X1_LVT execution_unit_0i_41_81 (.A1(execution_unit_0_n_41_65),.A2(execution_unit_0_n_41_66),.A3(execution_unit_0_n_41_67),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_68));
	AOI21_X1_LVT execution_unit_0i_41_82 (.A(execution_unit_0_n_41_68),.B1(cpu_halt_st),.B2(dbg_mem_dout[13]),.ZN(execution_unit_0_n_41_69));
	INV_X1_LVT execution_unit_0i_41_83 (.A(execution_unit_0_n_41_69),.ZN(execution_unit_0_n_91));
	NAND2_X1_LVT execution_unit_0i_41_72 (.A1(execution_unit_0_n_74),.A2(inst_sext[12]),.ZN(execution_unit_0_n_41_60));
	INV_X1_LVT execution_unit_0i_34_26 (.A(eu_mdb_in[12]),.ZN(execution_unit_0_n_34_14));
	NOR2_X1_LVT execution_unit_0i_34_27 (.A1(execution_unit_0_n_34_9),.A2(execution_unit_0_n_34_14),.ZN(execution_unit_0_n_62));
	NAND2_X1_LVT execution_unit_0i_41_73 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_62),.ZN(execution_unit_0_n_41_61));
	NAND2_X1_LVT execution_unit_0i_41_74 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[12]),.ZN(execution_unit_0_n_41_62));
	NAND4_X1_LVT execution_unit_0i_41_75 (.A1(execution_unit_0_n_41_60),.A2(execution_unit_0_n_41_61),.A3(execution_unit_0_n_41_62),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_63));
	AOI21_X1_LVT execution_unit_0i_41_76 (.A(execution_unit_0_n_41_63),.B1(cpu_halt_st),.B2(dbg_mem_dout[12]),.ZN(execution_unit_0_n_41_64));
	INV_X1_LVT execution_unit_0i_41_77 (.A(execution_unit_0_n_41_64),.ZN(execution_unit_0_n_90));
	NAND2_X1_LVT execution_unit_0i_41_66 (.A1(execution_unit_0_n_74),.A2(inst_sext[11]),.ZN(execution_unit_0_n_41_55));
	INV_X1_LVT execution_unit_0i_34_24 (.A(eu_mdb_in[11]),.ZN(execution_unit_0_n_34_13));
	NOR2_X1_LVT execution_unit_0i_34_25 (.A1(execution_unit_0_n_34_9),.A2(execution_unit_0_n_34_13),.ZN(execution_unit_0_n_61));
	NAND2_X1_LVT execution_unit_0i_41_67 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_61),.ZN(execution_unit_0_n_41_56));
	NAND2_X1_LVT execution_unit_0i_41_68 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[11]),.ZN(execution_unit_0_n_41_57));
	NAND4_X1_LVT execution_unit_0i_41_69 (.A1(execution_unit_0_n_41_55),.A2(execution_unit_0_n_41_56),.A3(execution_unit_0_n_41_57),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_58));
	AOI21_X1_LVT execution_unit_0i_41_70 (.A(execution_unit_0_n_41_58),.B1(cpu_halt_st),.B2(dbg_mem_dout[11]),.ZN(execution_unit_0_n_41_59));
	INV_X1_LVT execution_unit_0i_41_71 (.A(execution_unit_0_n_41_59),.ZN(execution_unit_0_n_89));
	NAND2_X1_LVT execution_unit_0i_41_60 (.A1(execution_unit_0_n_74),.A2(inst_sext[10]),.ZN(execution_unit_0_n_41_50));
	INV_X1_LVT execution_unit_0i_34_22 (.A(eu_mdb_in[10]),.ZN(execution_unit_0_n_34_12));
	NOR2_X1_LVT execution_unit_0i_34_23 (.A1(execution_unit_0_n_34_9),.A2(execution_unit_0_n_34_12),.ZN(execution_unit_0_n_60));
	NAND2_X1_LVT execution_unit_0i_41_61 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_60),.ZN(execution_unit_0_n_41_51));
	NAND2_X1_LVT execution_unit_0i_41_62 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[10]),.ZN(execution_unit_0_n_41_52));
	NAND4_X1_LVT execution_unit_0i_41_63 (.A1(execution_unit_0_n_41_50),.A2(execution_unit_0_n_41_51),.A3(execution_unit_0_n_41_52),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_53));
	AOI21_X1_LVT execution_unit_0i_41_64 (.A(execution_unit_0_n_41_53),.B1(cpu_halt_st),.B2(dbg_mem_dout[10]),.ZN(execution_unit_0_n_41_54));
	INV_X1_LVT execution_unit_0i_41_65 (.A(execution_unit_0_n_41_54),.ZN(execution_unit_0_n_88));
	NAND2_X1_LVT execution_unit_0i_41_54 (.A1(execution_unit_0_n_74),.A2(inst_sext[9]),.ZN(execution_unit_0_n_41_45));
	INV_X1_LVT execution_unit_0i_34_20 (.A(eu_mdb_in[9]),.ZN(execution_unit_0_n_34_11));
	NOR2_X1_LVT execution_unit_0i_34_21 (.A1(execution_unit_0_n_34_9),.A2(execution_unit_0_n_34_11),.ZN(execution_unit_0_n_59));
	NAND2_X1_LVT execution_unit_0i_41_55 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_59),.ZN(execution_unit_0_n_41_46));
	NAND2_X1_LVT execution_unit_0i_41_56 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[9]),.ZN(execution_unit_0_n_41_47));
	NAND4_X1_LVT execution_unit_0i_41_57 (.A1(execution_unit_0_n_41_45),.A2(execution_unit_0_n_41_46),.A3(execution_unit_0_n_41_47),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_48));
	AOI21_X1_LVT execution_unit_0i_41_58 (.A(execution_unit_0_n_41_48),.B1(cpu_halt_st),.B2(dbg_mem_dout[9]),.ZN(execution_unit_0_n_41_49));
	INV_X1_LVT execution_unit_0i_41_59 (.A(execution_unit_0_n_41_49),.ZN(execution_unit_0_n_87));
	NAND2_X1_LVT execution_unit_0i_41_48 (.A1(execution_unit_0_n_74),.A2(inst_sext[8]),.ZN(execution_unit_0_n_41_40));
	INV_X1_LVT execution_unit_0i_34_18 (.A(eu_mdb_in[8]),.ZN(execution_unit_0_n_34_10));
	NOR2_X1_LVT execution_unit_0i_34_19 (.A1(execution_unit_0_n_34_9),.A2(execution_unit_0_n_34_10),.ZN(execution_unit_0_n_58));
	NAND2_X1_LVT execution_unit_0i_41_49 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_58),.ZN(execution_unit_0_n_41_41));
	NAND2_X1_LVT execution_unit_0i_41_50 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[8]),.ZN(execution_unit_0_n_41_42));
	NAND4_X1_LVT execution_unit_0i_41_51 (.A1(execution_unit_0_n_41_40),.A2(execution_unit_0_n_41_41),.A3(execution_unit_0_n_41_42),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_43));
	AOI21_X1_LVT execution_unit_0i_41_52 (.A(execution_unit_0_n_41_43),.B1(cpu_halt_st),.B2(dbg_mem_dout[8]),.ZN(execution_unit_0_n_41_44));
	INV_X1_LVT execution_unit_0i_41_53 (.A(execution_unit_0_n_41_44),.ZN(execution_unit_0_n_86));
	NAND2_X1_LVT execution_unit_0i_41_42 (.A1(execution_unit_0_n_74),.A2(inst_sext[7]),.ZN(execution_unit_0_n_41_35));
	OR2_X1_LVT execution_unit_0i_34_0 (.A1(execution_unit_0_n_47),.A2(execution_unit_0_n_48),.ZN(execution_unit_0_n_34_0));
	AOI22_X1_LVT execution_unit_0i_34_15 (.A1(execution_unit_0_n_34_0),.A2(eu_mdb_in[7]),.B1(execution_unit_0_n_49),.B2(eu_mdb_in[15]),.ZN(execution_unit_0_n_34_8));
	INV_X1_LVT execution_unit_0i_34_16 (.A(execution_unit_0_n_34_8),.ZN(execution_unit_0_n_57));
	NAND2_X1_LVT execution_unit_0i_41_43 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_57),.ZN(execution_unit_0_n_41_36));
	NAND2_X1_LVT execution_unit_0i_41_44 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[7]),.ZN(execution_unit_0_n_41_37));
	NAND4_X1_LVT execution_unit_0i_41_45 (.A1(execution_unit_0_n_41_35),.A2(execution_unit_0_n_41_36),.A3(execution_unit_0_n_41_37),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_38));
	AOI21_X1_LVT execution_unit_0i_41_46 (.A(execution_unit_0_n_41_38),.B1(cpu_halt_st),.B2(dbg_mem_dout[7]),.ZN(execution_unit_0_n_41_39));
	INV_X1_LVT execution_unit_0i_41_47 (.A(execution_unit_0_n_41_39),.ZN(execution_unit_0_n_85));
	NAND2_X1_LVT execution_unit_0i_41_36 (.A1(execution_unit_0_n_74),.A2(inst_sext[6]),.ZN(execution_unit_0_n_41_30));
	AOI22_X1_LVT execution_unit_0i_34_13 (.A1(execution_unit_0_n_34_0),.A2(eu_mdb_in[6]),.B1(execution_unit_0_n_49),.B2(eu_mdb_in[14]),.ZN(execution_unit_0_n_34_7));
	INV_X1_LVT execution_unit_0i_34_14 (.A(execution_unit_0_n_34_7),.ZN(execution_unit_0_n_56));
	NAND2_X1_LVT execution_unit_0i_41_37 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_56),.ZN(execution_unit_0_n_41_31));
	NAND2_X1_LVT execution_unit_0i_41_38 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[6]),.ZN(execution_unit_0_n_41_32));
	NAND4_X1_LVT execution_unit_0i_41_39 (.A1(execution_unit_0_n_41_30),.A2(execution_unit_0_n_41_31),.A3(execution_unit_0_n_41_32),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_33));
	AOI21_X1_LVT execution_unit_0i_41_40 (.A(execution_unit_0_n_41_33),.B1(cpu_halt_st),.B2(dbg_mem_dout[6]),.ZN(execution_unit_0_n_41_34));
	INV_X1_LVT execution_unit_0i_41_41 (.A(execution_unit_0_n_41_34),.ZN(execution_unit_0_n_84));
	NAND2_X1_LVT execution_unit_0i_41_30 (.A1(execution_unit_0_n_74),.A2(inst_sext[5]),.ZN(execution_unit_0_n_41_25));
	AOI22_X1_LVT execution_unit_0i_34_11 (.A1(execution_unit_0_n_34_0),.A2(eu_mdb_in[5]),.B1(execution_unit_0_n_49),.B2(eu_mdb_in[13]),.ZN(execution_unit_0_n_34_6));
	INV_X1_LVT execution_unit_0i_34_12 (.A(execution_unit_0_n_34_6),.ZN(execution_unit_0_n_55));
	NAND2_X1_LVT execution_unit_0i_41_31 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_55),.ZN(execution_unit_0_n_41_26));
	NAND2_X1_LVT execution_unit_0i_41_32 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[5]),.ZN(execution_unit_0_n_41_27));
	NAND4_X1_LVT execution_unit_0i_41_33 (.A1(execution_unit_0_n_41_25),.A2(execution_unit_0_n_41_26),.A3(execution_unit_0_n_41_27),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_28));
	AOI21_X1_LVT execution_unit_0i_41_34 (.A(execution_unit_0_n_41_28),.B1(cpu_halt_st),.B2(dbg_mem_dout[5]),.ZN(execution_unit_0_n_41_29));
	INV_X1_LVT execution_unit_0i_41_35 (.A(execution_unit_0_n_41_29),.ZN(execution_unit_0_n_83));
	NAND2_X1_LVT execution_unit_0i_41_24 (.A1(execution_unit_0_n_74),.A2(inst_sext[4]),.ZN(execution_unit_0_n_41_20));
	AOI22_X1_LVT execution_unit_0i_34_9 (.A1(execution_unit_0_n_34_0),.A2(eu_mdb_in[4]),.B1(execution_unit_0_n_49),.B2(eu_mdb_in[12]),.ZN(execution_unit_0_n_34_5));
	INV_X1_LVT execution_unit_0i_34_10 (.A(execution_unit_0_n_34_5),.ZN(execution_unit_0_n_54));
	NAND2_X1_LVT execution_unit_0i_41_25 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_54),.ZN(execution_unit_0_n_41_21));
	NAND2_X1_LVT execution_unit_0i_41_26 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[4]),.ZN(execution_unit_0_n_41_22));
	NAND4_X1_LVT execution_unit_0i_41_27 (.A1(execution_unit_0_n_41_20),.A2(execution_unit_0_n_41_21),.A3(execution_unit_0_n_41_22),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_23));
	AOI21_X1_LVT execution_unit_0i_41_28 (.A(execution_unit_0_n_41_23),.B1(cpu_halt_st),.B2(dbg_mem_dout[4]),.ZN(execution_unit_0_n_41_24));
	INV_X1_LVT execution_unit_0i_41_29 (.A(execution_unit_0_n_41_24),.ZN(execution_unit_0_n_82));
	NAND2_X1_LVT execution_unit_0i_41_18 (.A1(execution_unit_0_n_74),.A2(inst_sext[3]),.ZN(execution_unit_0_n_41_15));
	AOI22_X1_LVT execution_unit_0i_34_7 (.A1(execution_unit_0_n_34_0),.A2(eu_mdb_in[3]),.B1(execution_unit_0_n_49),.B2(eu_mdb_in[11]),.ZN(execution_unit_0_n_34_4));
	INV_X1_LVT execution_unit_0i_34_8 (.A(execution_unit_0_n_34_4),.ZN(execution_unit_0_n_53));
	NAND2_X1_LVT execution_unit_0i_41_19 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_53),.ZN(execution_unit_0_n_41_16));
	NAND2_X1_LVT execution_unit_0i_41_20 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[3]),.ZN(execution_unit_0_n_41_17));
	NAND4_X1_LVT execution_unit_0i_41_21 (.A1(execution_unit_0_n_41_15),.A2(execution_unit_0_n_41_16),.A3(execution_unit_0_n_41_17),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_18));
	AOI21_X1_LVT execution_unit_0i_41_22 (.A(execution_unit_0_n_41_18),.B1(cpu_halt_st),.B2(dbg_mem_dout[3]),.ZN(execution_unit_0_n_41_19));
	INV_X1_LVT execution_unit_0i_41_23 (.A(execution_unit_0_n_41_19),.ZN(execution_unit_0_n_81));
	NAND2_X1_LVT execution_unit_0i_41_12 (.A1(execution_unit_0_n_74),.A2(inst_sext[2]),.ZN(execution_unit_0_n_41_10));
	AOI22_X1_LVT execution_unit_0i_34_5 (.A1(execution_unit_0_n_34_0),.A2(eu_mdb_in[2]),.B1(execution_unit_0_n_49),.B2(eu_mdb_in[10]),.ZN(execution_unit_0_n_34_3));
	INV_X1_LVT execution_unit_0i_34_6 (.A(execution_unit_0_n_34_3),.ZN(execution_unit_0_n_52));
	NAND2_X1_LVT execution_unit_0i_41_13 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_52),.ZN(execution_unit_0_n_41_11));
	NAND2_X1_LVT execution_unit_0i_41_14 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[2]),.ZN(execution_unit_0_n_41_12));
	NAND4_X1_LVT execution_unit_0i_41_15 (.A1(execution_unit_0_n_41_10),.A2(execution_unit_0_n_41_11),.A3(execution_unit_0_n_41_12),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_13));
	AOI21_X1_LVT execution_unit_0i_41_16 (.A(execution_unit_0_n_41_13),.B1(cpu_halt_st),.B2(dbg_mem_dout[2]),.ZN(execution_unit_0_n_41_14));
	INV_X1_LVT execution_unit_0i_41_17 (.A(execution_unit_0_n_41_14),.ZN(execution_unit_0_n_80));
	NAND2_X1_LVT execution_unit_0i_41_5 (.A1(execution_unit_0_n_74),.A2(inst_sext[1]),.ZN(execution_unit_0_n_41_4));
	AOI22_X1_LVT execution_unit_0i_34_3 (.A1(execution_unit_0_n_34_0),.A2(eu_mdb_in[1]),.B1(execution_unit_0_n_49),.B2(eu_mdb_in[9]),.ZN(execution_unit_0_n_34_2));
	INV_X1_LVT execution_unit_0i_34_4 (.A(execution_unit_0_n_34_2),.ZN(execution_unit_0_n_51));
	NAND2_X1_LVT execution_unit_0i_41_6 (.A1(execution_unit_0_n_75),.A2(execution_unit_0_n_51),.ZN(execution_unit_0_n_41_5));
	NAND2_X1_LVT execution_unit_0i_41_7 (.A1(execution_unit_0_n_76),.A2(dbg_reg_din[1]),.ZN(execution_unit_0_n_41_6));
	NAND4_X1_LVT execution_unit_0i_41_9 (.A1(execution_unit_0_n_41_4),.A2(execution_unit_0_n_41_5),.A3(execution_unit_0_n_41_6),.A4(execution_unit_0_n_41_7),.ZN(execution_unit_0_n_41_8));
	AOI21_X1_LVT execution_unit_0i_41_10 (.A(execution_unit_0_n_41_8),.B1(cpu_halt_st),.B2(dbg_mem_dout[1]),.ZN(execution_unit_0_n_41_9));
	INV_X1_LVT execution_unit_0i_41_11 (.A(execution_unit_0_n_41_9),.ZN(execution_unit_0_n_79));
	NAND2_X1_LVT execution_unit_0i_41_0 (.A1(dbg_mem_dout[0]),.A2(cpu_halt_st),.ZN(execution_unit_0_n_41_0));
	NAND2_X1_LVT execution_unit_0i_41_1 (.A1(inst_sext[0]),.A2(execution_unit_0_n_74),.ZN(execution_unit_0_n_41_1));
	AOI22_X1_LVT execution_unit_0i_34_1 (.A1(execution_unit_0_n_34_0),.A2(eu_mdb_in[0]),.B1(eu_mdb_in[8]),.B2(execution_unit_0_n_49),.ZN(execution_unit_0_n_34_1));
	INV_X1_LVT execution_unit_0i_34_2 (.A(execution_unit_0_n_34_1),.ZN(execution_unit_0_n_50));
	NAND2_X1_LVT execution_unit_0i_41_2 (.A1(execution_unit_0_n_50),.A2(execution_unit_0_n_75),.ZN(execution_unit_0_n_41_2));
	NAND2_X1_LVT execution_unit_0i_41_3 (.A1(dbg_reg_din[0]),.A2(execution_unit_0_n_76),.ZN(execution_unit_0_n_41_3));
	NAND4_X1_LVT execution_unit_0i_41_4 (.A1(execution_unit_0_n_41_0),.A2(execution_unit_0_n_41_1),.A3(execution_unit_0_n_41_2),.A4(execution_unit_0_n_41_3),.ZN(execution_unit_0_n_78));
	OR2_X1_LVT execution_unit_0i_48_8 (.A1(execution_unit_0_n_45),.A2(execution_unit_0_n_66),.ZN(execution_unit_0_n_102));
	NOR4_X1_LVT execution_unit_0i_0_13 (.A1(e_state[0]),.A2(e_state[1]),.A3(e_state[2]),.A4(e_state[3]),.ZN(execution_unit_0_reg_sr_clr));
	NOR2_X1_LVT execution_unit_0i_48_9 (.A1(execution_unit_0_reg_sr_clr),.A2(execution_unit_0_n_7),.ZN(execution_unit_0_n_48_5));
	INV_X1_LVT execution_unit_0i_48_10 (.A(inst_type[1]),.ZN(execution_unit_0_n_48_6));
	NAND3_X1_LVT execution_unit_0i_48_11 (.A1(execution_unit_0_n_48_6),.A2(inst_as[0]),.A3(execution_unit_0_n_0),.ZN(execution_unit_0_n_48_7));
	INV_X1_LVT execution_unit_0i_47_0 (.A(inst_as[6]),.ZN(execution_unit_0_n_98));
	NAND2_X1_LVT execution_unit_0i_48_12 (.A1(execution_unit_0_n_2),.A2(execution_unit_0_n_98),.ZN(execution_unit_0_n_48_8));
	NAND2_X1_LVT execution_unit_0i_48_13 (.A1(execution_unit_0_n_98),.A2(execution_unit_0_n_1),.ZN(execution_unit_0_n_48_9));
	NAND4_X1_LVT execution_unit_0i_48_14 (.A1(execution_unit_0_n_48_5),.A2(execution_unit_0_n_48_7),.A3(execution_unit_0_n_48_8),.A4(execution_unit_0_n_48_9),.ZN(execution_unit_0_n_103));
	NOR2_X1_LVT execution_unit_0i_49_0 (.A1(execution_unit_0_n_102),.A2(execution_unit_0_n_103),.ZN(execution_unit_0_n_49_0));
	INV_X1_LVT execution_unit_0i_49_8 (.A(execution_unit_0_n_49_0),.ZN(execution_unit_0_n_49_7));
	INV_X1_LVT execution_unit_0i_44_0 (.A(e_state[2]),.ZN(execution_unit_0_n_44_0));
	NAND4_X1_LVT execution_unit_0i_44_1 (.A1(execution_unit_0_n_44_0),.A2(e_state[0]),.A3(e_state[1]),.A4(e_state[3]),.ZN(execution_unit_0_n_44_1));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_en_reg (.D(execution_unit_0_n_1),.RN(execution_unit_0_n_18),.CK(cpu_mclk),.Q(execution_unit_0_mdb_in_buf_en),.QN());
	AND2_X1_LVT execution_unit_0i_44_2 (.A1(execution_unit_0_n_44_1),.A2(execution_unit_0_mdb_in_buf_en),.ZN(execution_unit_0_n_96));
	INV_X1_LVT execution_unit_0i_45_0 (.A(e_state[2]),.ZN(execution_unit_0_n_45_0));
	NAND4_X1_LVT execution_unit_0i_45_1 (.A1(execution_unit_0_n_45_0),.A2(e_state[0]),.A3(e_state[1]),.A4(e_state[3]),.ZN(execution_unit_0_n_45_1));
	NAND2_X1_LVT execution_unit_0i_45_2 (.A1(execution_unit_0_n_45_1),.A2(execution_unit_0_mdb_in_buf_en),.ZN(execution_unit_0_n_45_2));
	NAND2_X1_LVT execution_unit_0i_45_3 (.A1(execution_unit_0_n_45_2),.A2(execution_unit_0_n_45_1),.ZN(execution_unit_0_n_97));
	CLKGATETST_X1_LVT execution_unit_0clk_gate_mdb_in_buf_valid_reg (.CK(cpu_mclk),.E(execution_unit_0_n_97),.SE(1'b0),.GCK(execution_unit_0_n_95));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_valid_reg (.D(execution_unit_0_n_96),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_95),.Q(execution_unit_0_mdb_in_buf_valid),.QN());
	OAI21_X1_LVT execution_unit_0i_48_5 (.A(execution_unit_0_n_0),.B1(execution_unit_0_n_41),.B2(execution_unit_0_n_69),.ZN(execution_unit_0_n_48_3));
	AND2_X1_LVT execution_unit_0i_31_0 (.A1(execution_unit_0_n_4),.A2(inst_so[6]),.ZN(execution_unit_0_reg_sr_wr));
	INV_X1_LVT execution_unit_0i_48_6 (.A(execution_unit_0_reg_sr_wr),.ZN(execution_unit_0_n_48_4));
	NAND2_X1_LVT execution_unit_0i_48_7 (.A1(execution_unit_0_n_48_3),.A2(execution_unit_0_n_48_4),.ZN(execution_unit_0_n_101));
	NAND2_X1_LVT execution_unit_0i_49_1 (.A1(execution_unit_0_mdb_in_buf_valid),.A2(execution_unit_0_n_101),.ZN(execution_unit_0_n_49_1));
	NOR2_X1_LVT execution_unit_0i_49_9 (.A1(execution_unit_0_n_49_7),.A2(execution_unit_0_n_49_1),.ZN(execution_unit_0_n_105));
	CLKGATETST_X1_LVT execution_unit_0clk_gate_mdb_in_buf_reg (.CK(cpu_mclk),.E(execution_unit_0_mdb_in_buf_en),.SE(1'b0),.GCK(execution_unit_0_n_94));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b15___05F05d (.D(execution_unit_0_n_65),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[15]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_105 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[15]),.ZN(execution_unit_0_n_50_90));
	NAND2_X1_LVT execution_unit_0i_49_2 (.A1(execution_unit_0_n_49_0),.A2(execution_unit_0_n_49_1),.ZN(execution_unit_0_n_49_2));
	INV_X1_LVT execution_unit_0i_49_10 (.A(execution_unit_0_n_101),.ZN(execution_unit_0_n_49_8));
	NOR2_X1_LVT execution_unit_0i_49_11 (.A1(execution_unit_0_n_49_2),.A2(execution_unit_0_n_49_8),.ZN(execution_unit_0_n_106));
	NAND2_X1_LVT execution_unit_0i_50_106 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_65),.ZN(execution_unit_0_n_50_91));
	NOR2_X1_LVT execution_unit_0i_49_3 (.A1(execution_unit_0_n_49_2),.A2(execution_unit_0_n_101),.ZN(execution_unit_0_n_49_3));
	INV_X1_LVT execution_unit_0i_20_0 (.A(execution_unit_0_n_38),.ZN(execution_unit_0_n_39));
	NAND2_X1_LVT execution_unit_0i_48_2 (.A1(execution_unit_0_n_3),.A2(execution_unit_0_n_39),.ZN(execution_unit_0_n_48_1));
	INV_X1_LVT execution_unit_0i_48_3 (.A(execution_unit_0_n_4),.ZN(execution_unit_0_n_48_2));
	OAI21_X1_LVT execution_unit_0i_48_4 (.A(execution_unit_0_n_48_1),.B1(execution_unit_0_n_48_2),.B2(execution_unit_0_n_37),.ZN(execution_unit_0_n_100));
	AND2_X1_LVT execution_unit_0i_49_12 (.A1(execution_unit_0_n_49_3),.A2(execution_unit_0_n_100),.ZN(execution_unit_0_n_107));
	NAND2_X1_LVT execution_unit_0i_50_107 (.A1(execution_unit_0_n_107),.A2(inst_dext[15]),.ZN(execution_unit_0_n_50_92));
	INV_X1_LVT execution_unit_0i_49_4 (.A(execution_unit_0_n_100),.ZN(execution_unit_0_n_49_4));
	NAND2_X1_LVT execution_unit_0i_49_5 (.A1(execution_unit_0_n_49_3),.A2(execution_unit_0_n_49_4),.ZN(execution_unit_0_n_49_5));
	OR4_X1_LVT execution_unit_0i_48_0 (.A1(inst_as[7]),.A2(inst_as[5]),.A3(inst_type[1]),.A4(inst_so[6]),.ZN(execution_unit_0_n_48_0));
	AND2_X1_LVT execution_unit_0i_48_1 (.A1(execution_unit_0_n_48_0),.A2(execution_unit_0_n_0),.ZN(execution_unit_0_n_99));
	INV_X1_LVT execution_unit_0i_49_13 (.A(execution_unit_0_n_99),.ZN(execution_unit_0_n_49_9));
	NOR2_X1_LVT execution_unit_0i_49_14 (.A1(execution_unit_0_n_49_5),.A2(execution_unit_0_n_49_9),.ZN(execution_unit_0_n_108));
	NAND2_X1_LVT execution_unit_0i_50_108 (.A1(execution_unit_0_n_108),.A2(inst_sext[15]),.ZN(execution_unit_0_n_50_93));
	NAND4_X1_LVT execution_unit_0i_50_109 (.A1(execution_unit_0_n_50_90),.A2(execution_unit_0_n_50_91),.A3(execution_unit_0_n_50_92),.A4(execution_unit_0_n_50_93),.ZN(execution_unit_0_n_50_94));
	INV_X1_LVT execution_unit_0i_49_6 (.A(execution_unit_0_n_102),.ZN(execution_unit_0_n_49_6));
	NOR2_X1_LVT execution_unit_0i_49_7 (.A1(execution_unit_0_n_49_6),.A2(execution_unit_0_n_103),.ZN(execution_unit_0_n_104));
	AOI221_X1_LVT execution_unit_0i_50_110 (.A(execution_unit_0_n_50_94),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[15]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[15]),.ZN(execution_unit_0_n_50_95));
	INV_X1_LVT execution_unit_0i_50_111 (.A(execution_unit_0_n_50_95),.ZN(execution_unit_0_n_124));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b14___05F05d (.D(execution_unit_0_n_64),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[14]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_98 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[14]),.ZN(execution_unit_0_n_50_84));
	NAND2_X1_LVT execution_unit_0i_50_99 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_64),.ZN(execution_unit_0_n_50_85));
	NAND2_X1_LVT execution_unit_0i_50_100 (.A1(execution_unit_0_n_107),.A2(inst_dext[14]),.ZN(execution_unit_0_n_50_86));
	NAND2_X1_LVT execution_unit_0i_50_101 (.A1(execution_unit_0_n_108),.A2(inst_sext[14]),.ZN(execution_unit_0_n_50_87));
	NAND4_X1_LVT execution_unit_0i_50_102 (.A1(execution_unit_0_n_50_84),.A2(execution_unit_0_n_50_85),.A3(execution_unit_0_n_50_86),.A4(execution_unit_0_n_50_87),.ZN(execution_unit_0_n_50_88));
	AOI221_X1_LVT execution_unit_0i_50_103 (.A(execution_unit_0_n_50_88),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[14]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[14]),.ZN(execution_unit_0_n_50_89));
	INV_X1_LVT execution_unit_0i_50_104 (.A(execution_unit_0_n_50_89),.ZN(execution_unit_0_n_123));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b13___05F05d (.D(execution_unit_0_n_63),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[13]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_91 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[13]),.ZN(execution_unit_0_n_50_78));
	NAND2_X1_LVT execution_unit_0i_50_92 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_63),.ZN(execution_unit_0_n_50_79));
	NAND2_X1_LVT execution_unit_0i_50_93 (.A1(execution_unit_0_n_107),.A2(inst_dext[13]),.ZN(execution_unit_0_n_50_80));
	NAND2_X1_LVT execution_unit_0i_50_94 (.A1(execution_unit_0_n_108),.A2(inst_sext[13]),.ZN(execution_unit_0_n_50_81));
	NAND4_X1_LVT execution_unit_0i_50_95 (.A1(execution_unit_0_n_50_78),.A2(execution_unit_0_n_50_79),.A3(execution_unit_0_n_50_80),.A4(execution_unit_0_n_50_81),.ZN(execution_unit_0_n_50_82));
	AOI221_X1_LVT execution_unit_0i_50_96 (.A(execution_unit_0_n_50_82),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[13]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[13]),.ZN(execution_unit_0_n_50_83));
	INV_X1_LVT execution_unit_0i_50_97 (.A(execution_unit_0_n_50_83),.ZN(execution_unit_0_n_122));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b12___05F05d (.D(execution_unit_0_n_62),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[12]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_84 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[12]),.ZN(execution_unit_0_n_50_72));
	NAND2_X1_LVT execution_unit_0i_50_85 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_62),.ZN(execution_unit_0_n_50_73));
	NAND2_X1_LVT execution_unit_0i_50_86 (.A1(execution_unit_0_n_107),.A2(inst_dext[12]),.ZN(execution_unit_0_n_50_74));
	NAND2_X1_LVT execution_unit_0i_50_87 (.A1(execution_unit_0_n_108),.A2(inst_sext[12]),.ZN(execution_unit_0_n_50_75));
	NAND4_X1_LVT execution_unit_0i_50_88 (.A1(execution_unit_0_n_50_72),.A2(execution_unit_0_n_50_73),.A3(execution_unit_0_n_50_74),.A4(execution_unit_0_n_50_75),.ZN(execution_unit_0_n_50_76));
	AOI221_X1_LVT execution_unit_0i_50_89 (.A(execution_unit_0_n_50_76),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[12]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[12]),.ZN(execution_unit_0_n_50_77));
	INV_X1_LVT execution_unit_0i_50_90 (.A(execution_unit_0_n_50_77),.ZN(execution_unit_0_n_121));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b11___05F05d (.D(execution_unit_0_n_61),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[11]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_77 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[11]),.ZN(execution_unit_0_n_50_66));
	NAND2_X1_LVT execution_unit_0i_50_78 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_61),.ZN(execution_unit_0_n_50_67));
	NAND2_X1_LVT execution_unit_0i_50_79 (.A1(execution_unit_0_n_107),.A2(inst_dext[11]),.ZN(execution_unit_0_n_50_68));
	NAND2_X1_LVT execution_unit_0i_50_80 (.A1(execution_unit_0_n_108),.A2(inst_sext[11]),.ZN(execution_unit_0_n_50_69));
	NAND4_X1_LVT execution_unit_0i_50_81 (.A1(execution_unit_0_n_50_66),.A2(execution_unit_0_n_50_67),.A3(execution_unit_0_n_50_68),.A4(execution_unit_0_n_50_69),.ZN(execution_unit_0_n_50_70));
	AOI221_X1_LVT execution_unit_0i_50_82 (.A(execution_unit_0_n_50_70),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[11]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[11]),.ZN(execution_unit_0_n_50_71));
	INV_X1_LVT execution_unit_0i_50_83 (.A(execution_unit_0_n_50_71),.ZN(execution_unit_0_n_120));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b10___05F05d (.D(execution_unit_0_n_60),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[10]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_70 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[10]),.ZN(execution_unit_0_n_50_60));
	NAND2_X1_LVT execution_unit_0i_50_71 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_60),.ZN(execution_unit_0_n_50_61));
	NAND2_X1_LVT execution_unit_0i_50_72 (.A1(execution_unit_0_n_107),.A2(inst_dext[10]),.ZN(execution_unit_0_n_50_62));
	NAND2_X1_LVT execution_unit_0i_50_73 (.A1(execution_unit_0_n_108),.A2(inst_sext[10]),.ZN(execution_unit_0_n_50_63));
	NAND4_X1_LVT execution_unit_0i_50_74 (.A1(execution_unit_0_n_50_60),.A2(execution_unit_0_n_50_61),.A3(execution_unit_0_n_50_62),.A4(execution_unit_0_n_50_63),.ZN(execution_unit_0_n_50_64));
	AOI221_X1_LVT execution_unit_0i_50_75 (.A(execution_unit_0_n_50_64),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[10]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[10]),.ZN(execution_unit_0_n_50_65));
	INV_X1_LVT execution_unit_0i_50_76 (.A(execution_unit_0_n_50_65),.ZN(execution_unit_0_n_119));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b9___05F05d (.D(execution_unit_0_n_59),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[9]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_63 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[9]),.ZN(execution_unit_0_n_50_54));
	NAND2_X1_LVT execution_unit_0i_50_64 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_59),.ZN(execution_unit_0_n_50_55));
	NAND2_X1_LVT execution_unit_0i_50_65 (.A1(execution_unit_0_n_107),.A2(inst_dext[9]),.ZN(execution_unit_0_n_50_56));
	NAND2_X1_LVT execution_unit_0i_50_66 (.A1(execution_unit_0_n_108),.A2(inst_sext[9]),.ZN(execution_unit_0_n_50_57));
	NAND4_X1_LVT execution_unit_0i_50_67 (.A1(execution_unit_0_n_50_54),.A2(execution_unit_0_n_50_55),.A3(execution_unit_0_n_50_56),.A4(execution_unit_0_n_50_57),.ZN(execution_unit_0_n_50_58));
	AOI221_X1_LVT execution_unit_0i_50_68 (.A(execution_unit_0_n_50_58),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[9]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[9]),.ZN(execution_unit_0_n_50_59));
	INV_X1_LVT execution_unit_0i_50_69 (.A(execution_unit_0_n_50_59),.ZN(execution_unit_0_n_118));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b8___05F05d (.D(execution_unit_0_n_58),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[8]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_56 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[8]),.ZN(execution_unit_0_n_50_48));
	NAND2_X1_LVT execution_unit_0i_50_57 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_58),.ZN(execution_unit_0_n_50_49));
	NAND2_X1_LVT execution_unit_0i_50_58 (.A1(execution_unit_0_n_107),.A2(inst_dext[8]),.ZN(execution_unit_0_n_50_50));
	NAND2_X1_LVT execution_unit_0i_50_59 (.A1(execution_unit_0_n_108),.A2(inst_sext[8]),.ZN(execution_unit_0_n_50_51));
	NAND4_X1_LVT execution_unit_0i_50_60 (.A1(execution_unit_0_n_50_48),.A2(execution_unit_0_n_50_49),.A3(execution_unit_0_n_50_50),.A4(execution_unit_0_n_50_51),.ZN(execution_unit_0_n_50_52));
	AOI221_X1_LVT execution_unit_0i_50_61 (.A(execution_unit_0_n_50_52),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[8]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[8]),.ZN(execution_unit_0_n_50_53));
	INV_X1_LVT execution_unit_0i_50_62 (.A(execution_unit_0_n_50_53),.ZN(execution_unit_0_n_117));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b7___05F05d (.D(execution_unit_0_n_57),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[7]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_49 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[7]),.ZN(execution_unit_0_n_50_42));
	NAND2_X1_LVT execution_unit_0i_50_50 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_57),.ZN(execution_unit_0_n_50_43));
	NAND2_X1_LVT execution_unit_0i_50_51 (.A1(execution_unit_0_n_107),.A2(inst_dext[7]),.ZN(execution_unit_0_n_50_44));
	NAND2_X1_LVT execution_unit_0i_50_52 (.A1(execution_unit_0_n_108),.A2(inst_sext[7]),.ZN(execution_unit_0_n_50_45));
	NAND4_X1_LVT execution_unit_0i_50_53 (.A1(execution_unit_0_n_50_42),.A2(execution_unit_0_n_50_43),.A3(execution_unit_0_n_50_44),.A4(execution_unit_0_n_50_45),.ZN(execution_unit_0_n_50_46));
	AOI221_X1_LVT execution_unit_0i_50_54 (.A(execution_unit_0_n_50_46),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[7]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[7]),.ZN(execution_unit_0_n_50_47));
	INV_X1_LVT execution_unit_0i_50_55 (.A(execution_unit_0_n_50_47),.ZN(execution_unit_0_n_116));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b6___05F05d (.D(execution_unit_0_n_56),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[6]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_42 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[6]),.ZN(execution_unit_0_n_50_36));
	NAND2_X1_LVT execution_unit_0i_50_43 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_56),.ZN(execution_unit_0_n_50_37));
	NAND2_X1_LVT execution_unit_0i_50_44 (.A1(execution_unit_0_n_107),.A2(inst_dext[6]),.ZN(execution_unit_0_n_50_38));
	NAND2_X1_LVT execution_unit_0i_50_45 (.A1(execution_unit_0_n_108),.A2(inst_sext[6]),.ZN(execution_unit_0_n_50_39));
	NAND4_X1_LVT execution_unit_0i_50_46 (.A1(execution_unit_0_n_50_36),.A2(execution_unit_0_n_50_37),.A3(execution_unit_0_n_50_38),.A4(execution_unit_0_n_50_39),.ZN(execution_unit_0_n_50_40));
	AOI221_X1_LVT execution_unit_0i_50_47 (.A(execution_unit_0_n_50_40),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[6]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[6]),.ZN(execution_unit_0_n_50_41));
	INV_X1_LVT execution_unit_0i_50_48 (.A(execution_unit_0_n_50_41),.ZN(execution_unit_0_n_115));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b5___05F05d (.D(execution_unit_0_n_55),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[5]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_35 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[5]),.ZN(execution_unit_0_n_50_30));
	NAND2_X1_LVT execution_unit_0i_50_36 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_55),.ZN(execution_unit_0_n_50_31));
	NAND2_X1_LVT execution_unit_0i_50_37 (.A1(execution_unit_0_n_107),.A2(inst_dext[5]),.ZN(execution_unit_0_n_50_32));
	NAND2_X1_LVT execution_unit_0i_50_38 (.A1(execution_unit_0_n_108),.A2(inst_sext[5]),.ZN(execution_unit_0_n_50_33));
	NAND4_X1_LVT execution_unit_0i_50_39 (.A1(execution_unit_0_n_50_30),.A2(execution_unit_0_n_50_31),.A3(execution_unit_0_n_50_32),.A4(execution_unit_0_n_50_33),.ZN(execution_unit_0_n_50_34));
	AOI221_X1_LVT execution_unit_0i_50_40 (.A(execution_unit_0_n_50_34),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[5]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[5]),.ZN(execution_unit_0_n_50_35));
	INV_X1_LVT execution_unit_0i_50_41 (.A(execution_unit_0_n_50_35),.ZN(execution_unit_0_n_114));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b4___05F05d (.D(execution_unit_0_n_54),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[4]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_28 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[4]),.ZN(execution_unit_0_n_50_24));
	NAND2_X1_LVT execution_unit_0i_50_29 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_54),.ZN(execution_unit_0_n_50_25));
	NAND2_X1_LVT execution_unit_0i_50_30 (.A1(execution_unit_0_n_107),.A2(inst_dext[4]),.ZN(execution_unit_0_n_50_26));
	NAND2_X1_LVT execution_unit_0i_50_31 (.A1(execution_unit_0_n_108),.A2(inst_sext[4]),.ZN(execution_unit_0_n_50_27));
	NAND4_X1_LVT execution_unit_0i_50_32 (.A1(execution_unit_0_n_50_24),.A2(execution_unit_0_n_50_25),.A3(execution_unit_0_n_50_26),.A4(execution_unit_0_n_50_27),.ZN(execution_unit_0_n_50_28));
	AOI221_X1_LVT execution_unit_0i_50_33 (.A(execution_unit_0_n_50_28),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[4]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[4]),.ZN(execution_unit_0_n_50_29));
	INV_X1_LVT execution_unit_0i_50_34 (.A(execution_unit_0_n_50_29),.ZN(execution_unit_0_n_113));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b3___05F05d (.D(execution_unit_0_n_53),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[3]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_21 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[3]),.ZN(execution_unit_0_n_50_18));
	NAND2_X1_LVT execution_unit_0i_50_22 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_53),.ZN(execution_unit_0_n_50_19));
	NAND2_X1_LVT execution_unit_0i_50_23 (.A1(execution_unit_0_n_107),.A2(inst_dext[3]),.ZN(execution_unit_0_n_50_20));
	NAND2_X1_LVT execution_unit_0i_50_24 (.A1(execution_unit_0_n_108),.A2(inst_sext[3]),.ZN(execution_unit_0_n_50_21));
	NAND4_X1_LVT execution_unit_0i_50_25 (.A1(execution_unit_0_n_50_18),.A2(execution_unit_0_n_50_19),.A3(execution_unit_0_n_50_20),.A4(execution_unit_0_n_50_21),.ZN(execution_unit_0_n_50_22));
	AOI221_X1_LVT execution_unit_0i_50_26 (.A(execution_unit_0_n_50_22),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[3]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[3]),.ZN(execution_unit_0_n_50_23));
	INV_X1_LVT execution_unit_0i_50_27 (.A(execution_unit_0_n_50_23),.ZN(execution_unit_0_n_112));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b2___05F05d (.D(execution_unit_0_n_52),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[2]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_14 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[2]),.ZN(execution_unit_0_n_50_12));
	NAND2_X1_LVT execution_unit_0i_50_15 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_52),.ZN(execution_unit_0_n_50_13));
	NAND2_X1_LVT execution_unit_0i_50_16 (.A1(execution_unit_0_n_107),.A2(inst_dext[2]),.ZN(execution_unit_0_n_50_14));
	NAND2_X1_LVT execution_unit_0i_50_17 (.A1(execution_unit_0_n_108),.A2(inst_sext[2]),.ZN(execution_unit_0_n_50_15));
	NAND4_X1_LVT execution_unit_0i_50_18 (.A1(execution_unit_0_n_50_12),.A2(execution_unit_0_n_50_13),.A3(execution_unit_0_n_50_14),.A4(execution_unit_0_n_50_15),.ZN(execution_unit_0_n_50_16));
	AOI221_X1_LVT execution_unit_0i_50_19 (.A(execution_unit_0_n_50_16),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[2]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[2]),.ZN(execution_unit_0_n_50_17));
	INV_X1_LVT execution_unit_0i_50_20 (.A(execution_unit_0_n_50_17),.ZN(execution_unit_0_n_111));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b1___05F05d (.D(execution_unit_0_n_51),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[1]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_7 (.A1(execution_unit_0_n_105),.A2(execution_unit_0_mdb_in_buf[1]),.ZN(execution_unit_0_n_50_6));
	NAND2_X1_LVT execution_unit_0i_50_8 (.A1(execution_unit_0_n_106),.A2(execution_unit_0_n_51),.ZN(execution_unit_0_n_50_7));
	NAND2_X1_LVT execution_unit_0i_50_9 (.A1(execution_unit_0_n_107),.A2(inst_dext[1]),.ZN(execution_unit_0_n_50_8));
	NAND2_X1_LVT execution_unit_0i_50_10 (.A1(execution_unit_0_n_108),.A2(inst_sext[1]),.ZN(execution_unit_0_n_50_9));
	NAND4_X1_LVT execution_unit_0i_50_11 (.A1(execution_unit_0_n_50_6),.A2(execution_unit_0_n_50_7),.A3(execution_unit_0_n_50_8),.A4(execution_unit_0_n_50_9),.ZN(execution_unit_0_n_50_10));
	AOI221_X1_LVT execution_unit_0i_50_12 (.A(execution_unit_0_n_50_10),.B1(execution_unit_0_n_103),.B2(execution_unit_0_reg_src[1]),.C1(execution_unit_0_n_104),.C2(dbg_reg_din[1]),.ZN(execution_unit_0_n_50_11));
	INV_X1_LVT execution_unit_0i_50_13 (.A(execution_unit_0_n_50_11),.ZN(execution_unit_0_n_110));
	DFFR_X1_LVT execution_unit_0mdb_in_buf_reg___05F05b0___05F05d (.D(execution_unit_0_n_50),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_94),.Q(execution_unit_0_mdb_in_buf[0]),.QN());
	NAND2_X1_LVT execution_unit_0i_50_0 (.A1(execution_unit_0_mdb_in_buf[0]),.A2(execution_unit_0_n_105),.ZN(execution_unit_0_n_50_0));
	NAND2_X1_LVT execution_unit_0i_50_1 (.A1(execution_unit_0_n_50),.A2(execution_unit_0_n_106),.ZN(execution_unit_0_n_50_1));
	NAND2_X1_LVT execution_unit_0i_50_2 (.A1(inst_dext[0]),.A2(execution_unit_0_n_107),.ZN(execution_unit_0_n_50_2));
	NAND2_X1_LVT execution_unit_0i_50_3 (.A1(inst_sext[0]),.A2(execution_unit_0_n_108),.ZN(execution_unit_0_n_50_3));
	NAND4_X1_LVT execution_unit_0i_50_4 (.A1(execution_unit_0_n_50_0),.A2(execution_unit_0_n_50_1),.A3(execution_unit_0_n_50_2),.A4(execution_unit_0_n_50_3),.ZN(execution_unit_0_n_50_4));
	AOI221_X1_LVT execution_unit_0i_50_5 (.A(execution_unit_0_n_50_4),.B1(execution_unit_0_reg_src[0]),.B2(execution_unit_0_n_103),.C1(dbg_reg_din[0]),.C2(execution_unit_0_n_104),.ZN(execution_unit_0_n_50_5));
	INV_X1_LVT execution_unit_0i_50_6 (.A(execution_unit_0_n_50_5),.ZN(execution_unit_0_n_109));
	OR3_X1_LVT execution_unit_0alu_0i_42_0 (.A1(inst_so[7]),.A2(inst_alu[3]),.A3(cpu_halt_st),.ZN(execution_unit_0_alu_0_n_104));
	NAND2_X1_LVT execution_unit_0alu_0i_0_0 (.A1(execution_unit_0_n_0),.A2(inst_bw),.ZN(execution_unit_0_alu_0_op_bit8_msk));
	AND2_X1_LVT execution_unit_0alu_0i_1_7 (.A1(execution_unit_0_alu_0_op_bit8_msk),.A2(execution_unit_0_n_78),.ZN(execution_unit_0_alu_0_n_7));
	XOR2_X1_LVT execution_unit_0alu_0i_29_0 (.A(execution_unit_0_status[3]),.B(execution_unit_0_status[2]),.Z(execution_unit_0_alu_0_n_86));
	INV_X1_LVT execution_unit_0alu_0i_30_0 (.A(execution_unit_0_alu_0_n_86),.ZN(execution_unit_0_alu_0_n_30_0));
	INV_X1_LVT execution_unit_0alu_0i_30_1 (.A(execution_unit_0_status[1]),.ZN(execution_unit_0_alu_0_n_30_1));
	INV_X1_LVT execution_unit_0alu_0i_30_2 (.A(execution_unit_0_status[0]),.ZN(execution_unit_0_alu_0_n_30_2));
	AOI222_X1_LVT execution_unit_0alu_0i_30_3 (.A1(execution_unit_0_alu_0_n_30_0),.A2(inst_jmp[6]),.B1(execution_unit_0_alu_0_n_30_1),.B2(inst_jmp[1]),.C1(execution_unit_0_alu_0_n_30_2),.C2(inst_jmp[3]),.ZN(execution_unit_0_alu_0_n_30_3));
	INV_X1_LVT execution_unit_0alu_0i_30_4 (.A(execution_unit_0_status[2]),.ZN(execution_unit_0_alu_0_n_30_4));
	NAND2_X1_LVT execution_unit_0alu_0i_30_5 (.A1(execution_unit_0_alu_0_n_30_4),.A2(inst_jmp[4]),.ZN(execution_unit_0_alu_0_n_30_5));
	NAND2_X1_LVT execution_unit_0alu_0i_30_6 (.A1(inst_jmp[0]),.A2(execution_unit_0_status[1]),.ZN(execution_unit_0_alu_0_n_30_6));
	NAND2_X1_LVT execution_unit_0alu_0i_30_7 (.A1(inst_jmp[2]),.A2(execution_unit_0_status[0]),.ZN(execution_unit_0_alu_0_n_30_7));
	NAND2_X1_LVT execution_unit_0alu_0i_30_8 (.A1(execution_unit_0_alu_0_n_86),.A2(inst_jmp[5]),.ZN(execution_unit_0_alu_0_n_30_8));
	AND4_X1_LVT execution_unit_0alu_0i_30_9 (.A1(execution_unit_0_alu_0_n_30_5),.A2(execution_unit_0_alu_0_n_30_6),.A3(execution_unit_0_alu_0_n_30_7),.A4(execution_unit_0_alu_0_n_30_8),.ZN(execution_unit_0_alu_0_n_30_9));
	AND2_X1_LVT execution_unit_0alu_0i_30_10 (.A1(execution_unit_0_alu_0_n_30_3),.A2(execution_unit_0_alu_0_n_30_9),.ZN(execution_unit_0_alu_0_n_87));
	AND2_X1_LVT execution_unit_0alu_0i_2_0 (.A1(execution_unit_0_n_0),.A2(inst_alu[0]),.ZN(execution_unit_0_alu_0_op_src_inv_cmd));
	XNOR2_X1_LVT execution_unit_0alu_0i_4_15 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_109),.ZN(execution_unit_0_alu_0_n_4_8));
	INV_X1_LVT execution_unit_0alu_0i_4_1 (.A(execution_unit_0_alu_0_op_bit8_msk),.ZN(execution_unit_0_alu_0_n_4_1));
	NOR2_X1_LVT execution_unit_0alu_0i_4_16 (.A1(execution_unit_0_alu_0_n_4_8),.A2(execution_unit_0_alu_0_n_4_1),.ZN(execution_unit_0_alu_0_X[3]));
	AND2_X1_LVT execution_unit_0alu_0i_39_7 (.A1(execution_unit_0_alu_0_n_87),.A2(execution_unit_0_alu_0_X[3]),.ZN(execution_unit_0_alu_0_n_103));
	AND2_X1_LVT execution_unit_0alu_0i_1_6 (.A1(execution_unit_0_alu_0_op_bit8_msk),.A2(execution_unit_0_n_79),.ZN(execution_unit_0_alu_0_n_6));
	XNOR2_X1_LVT execution_unit_0alu_0i_4_13 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_110),.ZN(execution_unit_0_alu_0_n_4_7));
	NOR2_X1_LVT execution_unit_0alu_0i_4_14 (.A1(execution_unit_0_alu_0_n_4_7),.A2(execution_unit_0_alu_0_n_4_1),.ZN(execution_unit_0_alu_0_X[2]));
	AND2_X1_LVT execution_unit_0alu_0i_39_6 (.A1(execution_unit_0_alu_0_n_87),.A2(execution_unit_0_alu_0_X[2]),.ZN(execution_unit_0_alu_0_n_102));
	AND2_X1_LVT execution_unit_0alu_0i_1_5 (.A1(execution_unit_0_alu_0_op_bit8_msk),.A2(execution_unit_0_n_80),.ZN(execution_unit_0_alu_0_n_5));
	XNOR2_X1_LVT execution_unit_0alu_0i_4_11 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_111),.ZN(execution_unit_0_alu_0_n_4_6));
	NOR2_X1_LVT execution_unit_0alu_0i_4_12 (.A1(execution_unit_0_alu_0_n_4_6),.A2(execution_unit_0_alu_0_n_4_1),.ZN(execution_unit_0_alu_0_X[1]));
	AND2_X1_LVT execution_unit_0alu_0i_39_5 (.A1(execution_unit_0_alu_0_n_87),.A2(execution_unit_0_alu_0_X[1]),.ZN(execution_unit_0_alu_0_n_101));
	AND2_X1_LVT execution_unit_0alu_0i_1_4 (.A1(execution_unit_0_alu_0_op_bit8_msk),.A2(execution_unit_0_n_81),.ZN(execution_unit_0_alu_0_n_4));
	XNOR2_X1_LVT execution_unit_0alu_0i_4_9 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_112),.ZN(execution_unit_0_alu_0_n_4_5));
	NOR2_X1_LVT execution_unit_0alu_0i_4_10 (.A1(execution_unit_0_alu_0_n_4_5),.A2(execution_unit_0_alu_0_n_4_1),.ZN(execution_unit_0_alu_0_X[0]));
	AND2_X1_LVT execution_unit_0alu_0i_39_4 (.A1(execution_unit_0_alu_0_n_87),.A2(execution_unit_0_alu_0_X[0]),.ZN(execution_unit_0_alu_0_n_100));
	AND2_X1_LVT execution_unit_0alu_0i_1_3 (.A1(execution_unit_0_alu_0_op_bit8_msk),.A2(execution_unit_0_n_82),.ZN(execution_unit_0_alu_0_n_3));
	XNOR2_X1_LVT execution_unit_0alu_0i_4_7 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_113),.ZN(execution_unit_0_alu_0_n_4_4));
	NOR2_X1_LVT execution_unit_0alu_0i_4_8 (.A1(execution_unit_0_alu_0_n_4_4),.A2(execution_unit_0_alu_0_n_4_1),.ZN(execution_unit_0_alu_0_n_19));
	AND2_X1_LVT execution_unit_0alu_0i_39_3 (.A1(execution_unit_0_alu_0_n_87),.A2(execution_unit_0_alu_0_n_19),.ZN(execution_unit_0_alu_0_n_99));
	AND2_X1_LVT execution_unit_0alu_0i_1_2 (.A1(execution_unit_0_alu_0_op_bit8_msk),.A2(execution_unit_0_n_83),.ZN(execution_unit_0_alu_0_n_2));
	XNOR2_X1_LVT execution_unit_0alu_0i_4_5 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_114),.ZN(execution_unit_0_alu_0_n_4_3));
	NOR2_X1_LVT execution_unit_0alu_0i_4_6 (.A1(execution_unit_0_alu_0_n_4_3),.A2(execution_unit_0_alu_0_n_4_1),.ZN(execution_unit_0_alu_0_n_18));
	AND2_X1_LVT execution_unit_0alu_0i_39_2 (.A1(execution_unit_0_alu_0_n_87),.A2(execution_unit_0_alu_0_n_18),.ZN(execution_unit_0_alu_0_n_98));
	AND2_X1_LVT execution_unit_0alu_0i_1_1 (.A1(execution_unit_0_alu_0_op_bit8_msk),.A2(execution_unit_0_n_84),.ZN(execution_unit_0_alu_0_n_1));
	XNOR2_X1_LVT execution_unit_0alu_0i_4_3 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_115),.ZN(execution_unit_0_alu_0_n_4_2));
	NOR2_X1_LVT execution_unit_0alu_0i_4_4 (.A1(execution_unit_0_alu_0_n_4_2),.A2(execution_unit_0_alu_0_n_4_1),.ZN(execution_unit_0_alu_0_n_17));
	AND2_X1_LVT execution_unit_0alu_0i_39_1 (.A1(execution_unit_0_alu_0_n_87),.A2(execution_unit_0_alu_0_n_17),.ZN(execution_unit_0_alu_0_n_97));
	AND2_X1_LVT execution_unit_0alu_0i_1_0 (.A1(execution_unit_0_n_85),.A2(execution_unit_0_alu_0_op_bit8_msk),.ZN(execution_unit_0_alu_0_n_0));
	XNOR2_X1_LVT execution_unit_0alu_0i_4_0 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_116),.ZN(execution_unit_0_alu_0_n_4_0));
	NOR2_X1_LVT execution_unit_0alu_0i_4_2 (.A1(execution_unit_0_alu_0_n_4_0),.A2(execution_unit_0_alu_0_n_4_1),.ZN(execution_unit_0_alu_0_n_16));
	AND2_X1_LVT execution_unit_0alu_0i_39_0 (.A1(execution_unit_0_alu_0_n_16),.A2(execution_unit_0_alu_0_n_87),.ZN(execution_unit_0_alu_0_n_96));
	XOR2_X1_LVT execution_unit_0alu_0i_3_7 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_117),.Z(execution_unit_0_alu_0_n_15));
	AND2_X1_LVT execution_unit_0alu_0i_38_0 (.A1(execution_unit_0_alu_0_n_15),.A2(execution_unit_0_alu_0_n_87),.ZN(execution_unit_0_alu_0_n_95));
	XOR2_X1_LVT execution_unit_0alu_0i_3_6 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_118),.Z(execution_unit_0_alu_0_n_14));
	AND2_X1_LVT execution_unit_0alu_0i_37_0 (.A1(execution_unit_0_alu_0_n_14),.A2(execution_unit_0_alu_0_n_87),.ZN(execution_unit_0_alu_0_n_94));
	XOR2_X1_LVT execution_unit_0alu_0i_3_5 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_119),.Z(execution_unit_0_alu_0_n_13));
	AND2_X1_LVT execution_unit_0alu_0i_36_0 (.A1(execution_unit_0_alu_0_n_13),.A2(execution_unit_0_alu_0_n_87),.ZN(execution_unit_0_alu_0_n_93));
	XOR2_X1_LVT execution_unit_0alu_0i_3_4 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_120),.Z(execution_unit_0_alu_0_n_12));
	AND2_X1_LVT execution_unit_0alu_0i_35_0 (.A1(execution_unit_0_alu_0_n_12),.A2(execution_unit_0_alu_0_n_87),.ZN(execution_unit_0_alu_0_n_92));
	XOR2_X1_LVT execution_unit_0alu_0i_3_3 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_121),.Z(execution_unit_0_alu_0_n_11));
	AND2_X1_LVT execution_unit_0alu_0i_34_0 (.A1(execution_unit_0_alu_0_n_11),.A2(execution_unit_0_alu_0_n_87),.ZN(execution_unit_0_alu_0_n_91));
	XOR2_X1_LVT execution_unit_0alu_0i_3_2 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_122),.Z(execution_unit_0_alu_0_n_10));
	AND2_X1_LVT execution_unit_0alu_0i_33_0 (.A1(execution_unit_0_alu_0_n_10),.A2(execution_unit_0_alu_0_n_87),.ZN(execution_unit_0_alu_0_n_90));
	XOR2_X1_LVT execution_unit_0alu_0i_3_1 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_123),.Z(execution_unit_0_alu_0_n_9));
	AND2_X1_LVT execution_unit_0alu_0i_32_0 (.A1(execution_unit_0_alu_0_n_9),.A2(execution_unit_0_alu_0_n_87),.ZN(execution_unit_0_alu_0_n_89));
	XOR2_X1_LVT execution_unit_0alu_0i_3_0 (.A(execution_unit_0_alu_0_op_src_inv_cmd),.B(execution_unit_0_n_124),.Z(execution_unit_0_alu_0_n_8));
	AND2_X1_LVT execution_unit_0alu_0i_31_0 (.A1(execution_unit_0_alu_0_n_8),.A2(execution_unit_0_alu_0_n_87),.ZN(execution_unit_0_alu_0_n_88));
	HA_X1_LVT execution_unit_0alu_0i_40_0 (.A(execution_unit_0_n_93),.B(execution_unit_0_alu_0_n_88),.CO(execution_unit_0_alu_0_n_40_0),.S(eu_mab[0]));
	FA_X1_LVT execution_unit_0alu_0i_40_1 (.A(execution_unit_0_n_92),.B(execution_unit_0_alu_0_n_89),.CI(execution_unit_0_alu_0_n_40_0),.CO(execution_unit_0_alu_0_n_40_1),.S(eu_mab[1]));
	FA_X1_LVT execution_unit_0alu_0i_40_2 (.A(execution_unit_0_n_91),.B(execution_unit_0_alu_0_n_90),.CI(execution_unit_0_alu_0_n_40_1),.CO(execution_unit_0_alu_0_n_40_2),.S(eu_mab[2]));
	FA_X1_LVT execution_unit_0alu_0i_40_3 (.A(execution_unit_0_n_90),.B(execution_unit_0_alu_0_n_91),.CI(execution_unit_0_alu_0_n_40_2),.CO(execution_unit_0_alu_0_n_40_3),.S(eu_mab[3]));
	FA_X1_LVT execution_unit_0alu_0i_40_4 (.A(execution_unit_0_n_89),.B(execution_unit_0_alu_0_n_92),.CI(execution_unit_0_alu_0_n_40_3),.CO(execution_unit_0_alu_0_n_40_4),.S(eu_mab[4]));
	FA_X1_LVT execution_unit_0alu_0i_40_5 (.A(execution_unit_0_n_88),.B(execution_unit_0_alu_0_n_93),.CI(execution_unit_0_alu_0_n_40_4),.CO(execution_unit_0_alu_0_n_40_5),.S(eu_mab[5]));
	FA_X1_LVT execution_unit_0alu_0i_40_6 (.A(execution_unit_0_n_87),.B(execution_unit_0_alu_0_n_94),.CI(execution_unit_0_alu_0_n_40_5),.CO(execution_unit_0_alu_0_n_40_6),.S(eu_mab[6]));
	FA_X1_LVT execution_unit_0alu_0i_40_7 (.A(execution_unit_0_n_86),.B(execution_unit_0_alu_0_n_95),.CI(execution_unit_0_alu_0_n_40_6),.CO(execution_unit_0_alu_0_n_40_7),.S(eu_mab[7]));
	FA_X1_LVT execution_unit_0alu_0i_40_8 (.A(execution_unit_0_alu_0_n_0),.B(execution_unit_0_alu_0_n_96),.CI(execution_unit_0_alu_0_n_40_7),.CO(execution_unit_0_alu_0_n_40_8),.S(eu_mab[8]));
	FA_X1_LVT execution_unit_0alu_0i_40_9 (.A(execution_unit_0_alu_0_n_1),.B(execution_unit_0_alu_0_n_97),.CI(execution_unit_0_alu_0_n_40_8),.CO(execution_unit_0_alu_0_n_40_9),.S(eu_mab[9]));
	FA_X1_LVT execution_unit_0alu_0i_40_10 (.A(execution_unit_0_alu_0_n_2),.B(execution_unit_0_alu_0_n_98),.CI(execution_unit_0_alu_0_n_40_9),.CO(execution_unit_0_alu_0_n_40_10),.S(eu_mab[10]));
	FA_X1_LVT execution_unit_0alu_0i_40_11 (.A(execution_unit_0_alu_0_n_3),.B(execution_unit_0_alu_0_n_99),.CI(execution_unit_0_alu_0_n_40_10),.CO(execution_unit_0_alu_0_n_40_11),.S(eu_mab[11]));
	FA_X1_LVT execution_unit_0alu_0i_40_12 (.A(execution_unit_0_alu_0_n_4),.B(execution_unit_0_alu_0_n_100),.CI(execution_unit_0_alu_0_n_40_11),.CO(execution_unit_0_alu_0_n_40_12),.S(eu_mab[12]));
	FA_X1_LVT execution_unit_0alu_0i_40_13 (.A(execution_unit_0_alu_0_n_5),.B(execution_unit_0_alu_0_n_101),.CI(execution_unit_0_alu_0_n_40_12),.CO(execution_unit_0_alu_0_n_40_13),.S(eu_mab[13]));
	FA_X1_LVT execution_unit_0alu_0i_40_14 (.A(execution_unit_0_alu_0_n_6),.B(execution_unit_0_alu_0_n_102),.CI(execution_unit_0_alu_0_n_40_13),.CO(execution_unit_0_alu_0_n_40_14),.S(eu_mab[14]));
	FA_X1_LVT execution_unit_0alu_0i_40_15 (.A(execution_unit_0_alu_0_n_7),.B(execution_unit_0_alu_0_n_103),.CI(execution_unit_0_alu_0_n_40_14),.CO(execution_unit_0_alu_0_alu_add[0]),.S(eu_mab[15]));
	AOI21_X1_LVT execution_unit_0alu_0i_28_0 (.A(inst_alu[1]),.B1(inst_alu[2]),.B2(execution_unit_0_status[0]),.ZN(execution_unit_0_alu_0_n_28_0));
	INV_X1_LVT execution_unit_0alu_0i_28_1 (.A(execution_unit_0_n_0),.ZN(execution_unit_0_alu_0_n_28_1));
	NOR2_X1_LVT execution_unit_0alu_0i_28_2 (.A1(execution_unit_0_alu_0_n_28_0),.A2(execution_unit_0_alu_0_n_28_1),.ZN(execution_unit_0_alu_0_alu_inc));
	HA_X1_LVT execution_unit_0alu_0i_41_0 (.A(execution_unit_0_alu_0_alu_inc),.B(eu_mab[0]),.CO(execution_unit_0_alu_0_n_41_0),.S(execution_unit_0_alu_0_alu_add_inc[0]));
	HA_X1_LVT execution_unit_0alu_0i_41_1 (.A(eu_mab[1]),.B(execution_unit_0_alu_0_n_41_0),.CO(execution_unit_0_alu_0_n_41_1),.S(execution_unit_0_alu_0_alu_add_inc[1]));
	HA_X1_LVT execution_unit_0alu_0i_41_2 (.A(eu_mab[2]),.B(execution_unit_0_alu_0_n_41_1),.CO(execution_unit_0_alu_0_n_41_2),.S(execution_unit_0_alu_0_alu_add_inc[2]));
	HA_X1_LVT execution_unit_0alu_0i_41_3 (.A(eu_mab[3]),.B(execution_unit_0_alu_0_n_41_2),.CO(execution_unit_0_alu_0_n_41_3),.S(execution_unit_0_alu_0_alu_add_inc[3]));
	HA_X1_LVT execution_unit_0alu_0i_41_4 (.A(eu_mab[4]),.B(execution_unit_0_alu_0_n_41_3),.CO(execution_unit_0_alu_0_n_41_4),.S(execution_unit_0_alu_0_alu_add_inc[4]));
	HA_X1_LVT execution_unit_0alu_0i_41_5 (.A(eu_mab[5]),.B(execution_unit_0_alu_0_n_41_4),.CO(execution_unit_0_alu_0_n_41_5),.S(execution_unit_0_alu_0_alu_add_inc[5]));
	HA_X1_LVT execution_unit_0alu_0i_41_6 (.A(eu_mab[6]),.B(execution_unit_0_alu_0_n_41_5),.CO(execution_unit_0_alu_0_n_41_6),.S(execution_unit_0_alu_0_alu_add_inc[6]));
	HA_X1_LVT execution_unit_0alu_0i_41_7 (.A(eu_mab[7]),.B(execution_unit_0_alu_0_n_41_6),.CO(execution_unit_0_alu_0_n_41_7),.S(execution_unit_0_alu_0_alu_add_inc[7]));
	HA_X1_LVT execution_unit_0alu_0i_41_8 (.A(eu_mab[8]),.B(execution_unit_0_alu_0_n_41_7),.CO(execution_unit_0_alu_0_n_41_8),.S(execution_unit_0_alu_0_alu_add_inc[8]));
	HA_X1_LVT execution_unit_0alu_0i_41_9 (.A(eu_mab[9]),.B(execution_unit_0_alu_0_n_41_8),.CO(execution_unit_0_alu_0_n_41_9),.S(execution_unit_0_alu_0_alu_add_inc[9]));
	HA_X1_LVT execution_unit_0alu_0i_41_10 (.A(eu_mab[10]),.B(execution_unit_0_alu_0_n_41_9),.CO(execution_unit_0_alu_0_n_41_10),.S(execution_unit_0_alu_0_alu_add_inc[10]));
	HA_X1_LVT execution_unit_0alu_0i_41_11 (.A(eu_mab[11]),.B(execution_unit_0_alu_0_n_41_10),.CO(execution_unit_0_alu_0_n_41_11),.S(execution_unit_0_alu_0_alu_add_inc[11]));
	HA_X1_LVT execution_unit_0alu_0i_41_12 (.A(eu_mab[12]),.B(execution_unit_0_alu_0_n_41_11),.CO(execution_unit_0_alu_0_n_41_12),.S(execution_unit_0_alu_0_alu_add_inc[12]));
	HA_X1_LVT execution_unit_0alu_0i_41_13 (.A(eu_mab[13]),.B(execution_unit_0_alu_0_n_41_12),.CO(execution_unit_0_alu_0_n_41_13),.S(execution_unit_0_alu_0_alu_add_inc[13]));
	HA_X1_LVT execution_unit_0alu_0i_41_14 (.A(eu_mab[14]),.B(execution_unit_0_alu_0_n_41_13),.CO(execution_unit_0_alu_0_n_41_14),.S(execution_unit_0_alu_0_alu_add_inc[14]));
	HA_X1_LVT execution_unit_0alu_0i_41_15 (.A(eu_mab[15]),.B(execution_unit_0_alu_0_n_41_14),.CO(execution_unit_0_alu_0_n_41_15),.S(execution_unit_0_alu_0_alu_add_inc[15]));
	INV_X1_LVT execution_unit_0alu_0i_43_1 (.A(inst_alu[7]),.ZN(execution_unit_0_alu_0_n_43_0));
	NOR2_X1_LVT execution_unit_0alu_0i_43_2 (.A1(execution_unit_0_alu_0_n_43_0),.A2(execution_unit_0_alu_0_n_104),.ZN(execution_unit_0_alu_0_n_106));
	HA_X1_LVT execution_unit_0alu_0i_18_3 (.A(execution_unit_0_alu_0_n_3),.B(execution_unit_0_alu_0_n_19),.CO(execution_unit_0_alu_0_n_68),.S(execution_unit_0_alu_0_n_67));
	INV_X1_LVT execution_unit_0alu_0i_19_2 (.A(execution_unit_0_alu_0_n_68),.ZN(execution_unit_0_alu_0_n_19_3));
	HA_X1_LVT execution_unit_0alu_0i_18_2 (.A(execution_unit_0_alu_0_n_2),.B(execution_unit_0_alu_0_n_18),.CO(execution_unit_0_alu_0_n_66),.S(execution_unit_0_alu_0_n_65));
	HA_X1_LVT execution_unit_0alu_0i_19_1 (.A(execution_unit_0_alu_0_n_67),.B(execution_unit_0_alu_0_n_66),.CO(execution_unit_0_alu_0_n_19_2),.S(execution_unit_0_alu_0_n_19_1));
	HA_X1_LVT execution_unit_0alu_0i_13_3 (.A(execution_unit_0_n_86),.B(execution_unit_0_alu_0_n_15),.CO(execution_unit_0_alu_0_n_56),.S(execution_unit_0_alu_0_n_55));
	INV_X1_LVT execution_unit_0alu_0i_14_2 (.A(execution_unit_0_alu_0_n_56),.ZN(execution_unit_0_alu_0_n_14_3));
	HA_X1_LVT execution_unit_0alu_0i_13_2 (.A(execution_unit_0_n_87),.B(execution_unit_0_alu_0_n_14),.CO(execution_unit_0_alu_0_n_54),.S(execution_unit_0_alu_0_n_53));
	HA_X1_LVT execution_unit_0alu_0i_14_1 (.A(execution_unit_0_alu_0_n_55),.B(execution_unit_0_alu_0_n_54),.CO(execution_unit_0_alu_0_n_14_2),.S(execution_unit_0_alu_0_n_14_1));
	HA_X1_LVT execution_unit_0alu_0i_8_3 (.A(execution_unit_0_n_90),.B(execution_unit_0_alu_0_n_11),.CO(execution_unit_0_alu_0_n_44),.S(execution_unit_0_alu_0_n_43));
	INV_X1_LVT execution_unit_0alu_0i_9_2 (.A(execution_unit_0_alu_0_n_44),.ZN(execution_unit_0_alu_0_n_9_3));
	HA_X1_LVT execution_unit_0alu_0i_8_2 (.A(execution_unit_0_n_91),.B(execution_unit_0_alu_0_n_10),.CO(execution_unit_0_alu_0_n_42),.S(execution_unit_0_alu_0_n_41));
	HA_X1_LVT execution_unit_0alu_0i_9_1 (.A(execution_unit_0_alu_0_n_43),.B(execution_unit_0_alu_0_n_42),.CO(execution_unit_0_alu_0_n_9_2),.S(execution_unit_0_alu_0_n_9_1));
	FA_X1_LVT execution_unit_0alu_0i_8_0 (.A(execution_unit_0_n_93),.B(execution_unit_0_status[0]),.CI(execution_unit_0_alu_0_n_8),.CO(execution_unit_0_alu_0_n_8_0),.S(execution_unit_0_alu_0_n_38));
	FA_X1_LVT execution_unit_0alu_0i_8_1 (.A(execution_unit_0_n_92),.B(execution_unit_0_alu_0_n_9),.CI(execution_unit_0_alu_0_n_8_0),.CO(execution_unit_0_alu_0_n_40),.S(execution_unit_0_alu_0_n_39));
	INV_X1_LVT execution_unit_0alu_0i_9_0 (.A(execution_unit_0_alu_0_n_40),.ZN(execution_unit_0_alu_0_n_9_0));
	FA_X1_LVT execution_unit_0alu_0i_9_3 (.A(execution_unit_0_alu_0_n_41),.B(execution_unit_0_alu_0_n_9_0),.CI(execution_unit_0_alu_0_n_39),.CO(execution_unit_0_alu_0_n_9_4),.S());
	FA_X1_LVT execution_unit_0alu_0i_9_4 (.A(execution_unit_0_alu_0_n_40),.B(execution_unit_0_alu_0_n_9_1),.CI(execution_unit_0_alu_0_n_9_4),.CO(execution_unit_0_alu_0_n_9_5),.S());
	FA_X1_LVT execution_unit_0alu_0i_9_5 (.A(execution_unit_0_alu_0_n_9_2),.B(execution_unit_0_alu_0_n_9_3),.CI(execution_unit_0_alu_0_n_9_5),.CO(execution_unit_0_alu_0_n_9_6),.S());
	HA_X1_LVT execution_unit_0alu_0i_9_6 (.A(execution_unit_0_alu_0_n_9_3),.B(execution_unit_0_alu_0_n_9_6),.CO(execution_unit_0_alu_0_n_9_7),.S());
	HA_X1_LVT execution_unit_0alu_0i_9_7 (.A(execution_unit_0_alu_0_n_9_3),.B(execution_unit_0_alu_0_n_9_7),.CO(execution_unit_0_alu_0_n_9_8),.S());
	XNOR2_X1_LVT execution_unit_0alu_0i_9_8 (.A(execution_unit_0_alu_0_n_9_3),.B(execution_unit_0_alu_0_n_9_8),.ZN(execution_unit_0_alu_0_n_9_9));
	INV_X1_LVT execution_unit_0alu_0i_9_9 (.A(execution_unit_0_alu_0_n_9_9),.ZN(execution_unit_0_alu_0_n_45));
	INV_X1_LVT execution_unit_0alu_0i_10_0 (.A(execution_unit_0_alu_0_n_45),.ZN(execution_unit_0_alu_0_n_46));
	HA_X1_LVT execution_unit_0alu_0i_11_0 (.A(execution_unit_0_alu_0_n_40),.B(execution_unit_0_alu_0_n_41),.CO(execution_unit_0_alu_0_n_11_0),.S(execution_unit_0_alu_0_n_47));
	FA_X1_LVT execution_unit_0alu_0i_11_1 (.A(execution_unit_0_alu_0_n_43),.B(execution_unit_0_alu_0_n_42),.CI(execution_unit_0_alu_0_n_11_0),.CO(execution_unit_0_alu_0_n_11_1),.S(execution_unit_0_alu_0_n_48));
	OR2_X1_LVT execution_unit_0alu_0i_12_7 (.A1(execution_unit_0_alu_0_n_46),.A2(execution_unit_0_alu_0_n_48),.ZN(execution_unit_0_alu_0_n_12_5));
	HA_X1_LVT execution_unit_0alu_0i_11_2 (.A(execution_unit_0_alu_0_n_44),.B(execution_unit_0_alu_0_n_11_1),.CO(execution_unit_0_alu_0_n_11_2),.S(execution_unit_0_alu_0_n_49));
	INV_X1_LVT execution_unit_0alu_0i_12_8 (.A(execution_unit_0_alu_0_n_49),.ZN(execution_unit_0_alu_0_n_12_6));
	XNOR2_X1_LVT execution_unit_0alu_0i_12_10 (.A(execution_unit_0_alu_0_n_12_5),.B(execution_unit_0_alu_0_n_12_6),.ZN(execution_unit_0_alu_0_n_12_8));
	INV_X1_LVT execution_unit_0alu_0i_12_3 (.A(execution_unit_0_alu_0_n_39),.ZN(execution_unit_0_alu_0_n_12_2));
	NAND2_X1_LVT execution_unit_0alu_0i_12_2 (.A1(execution_unit_0_alu_0_n_46),.A2(execution_unit_0_alu_0_n_12_2),.ZN(execution_unit_0_alu_0_n_12_1));
	OR2_X1_LVT execution_unit_0alu_0i_12_5 (.A1(execution_unit_0_alu_0_n_47),.A2(execution_unit_0_alu_0_n_12_1),.ZN(execution_unit_0_alu_0_n_12_3));
	XNOR2_X1_LVT execution_unit_0alu_0i_12_6 (.A(execution_unit_0_alu_0_n_46),.B(execution_unit_0_alu_0_n_48),.ZN(execution_unit_0_alu_0_n_12_4));
	HA_X1_LVT execution_unit_0alu_0i_12_9 (.A(execution_unit_0_alu_0_n_12_3),.B(execution_unit_0_alu_0_n_12_4),.CO(execution_unit_0_alu_0_n_12_7),.S(execution_unit_0_alu_0_bcd_add[3]));
	XNOR2_X1_LVT execution_unit_0alu_0i_12_11 (.A(execution_unit_0_alu_0_n_12_8),.B(execution_unit_0_alu_0_n_12_7),.ZN(execution_unit_0_alu_0_bcd_add[4]));
	FA_X1_LVT execution_unit_0alu_0i_13_0 (.A(execution_unit_0_n_89),.B(execution_unit_0_alu_0_bcd_add[4]),.CI(execution_unit_0_alu_0_n_12),.CO(execution_unit_0_alu_0_n_13_0),.S(execution_unit_0_alu_0_n_50));
	FA_X1_LVT execution_unit_0alu_0i_13_1 (.A(execution_unit_0_n_88),.B(execution_unit_0_alu_0_n_13),.CI(execution_unit_0_alu_0_n_13_0),.CO(execution_unit_0_alu_0_n_52),.S(execution_unit_0_alu_0_n_51));
	INV_X1_LVT execution_unit_0alu_0i_14_0 (.A(execution_unit_0_alu_0_n_52),.ZN(execution_unit_0_alu_0_n_14_0));
	FA_X1_LVT execution_unit_0alu_0i_14_3 (.A(execution_unit_0_alu_0_n_53),.B(execution_unit_0_alu_0_n_14_0),.CI(execution_unit_0_alu_0_n_51),.CO(execution_unit_0_alu_0_n_14_4),.S());
	FA_X1_LVT execution_unit_0alu_0i_14_4 (.A(execution_unit_0_alu_0_n_52),.B(execution_unit_0_alu_0_n_14_1),.CI(execution_unit_0_alu_0_n_14_4),.CO(execution_unit_0_alu_0_n_14_5),.S());
	FA_X1_LVT execution_unit_0alu_0i_14_5 (.A(execution_unit_0_alu_0_n_14_2),.B(execution_unit_0_alu_0_n_14_3),.CI(execution_unit_0_alu_0_n_14_5),.CO(execution_unit_0_alu_0_n_14_6),.S());
	HA_X1_LVT execution_unit_0alu_0i_14_6 (.A(execution_unit_0_alu_0_n_14_3),.B(execution_unit_0_alu_0_n_14_6),.CO(execution_unit_0_alu_0_n_14_7),.S());
	HA_X1_LVT execution_unit_0alu_0i_14_7 (.A(execution_unit_0_alu_0_n_14_3),.B(execution_unit_0_alu_0_n_14_7),.CO(execution_unit_0_alu_0_n_14_8),.S());
	XNOR2_X1_LVT execution_unit_0alu_0i_14_8 (.A(execution_unit_0_alu_0_n_14_3),.B(execution_unit_0_alu_0_n_14_8),.ZN(execution_unit_0_alu_0_n_14_9));
	INV_X1_LVT execution_unit_0alu_0i_14_9 (.A(execution_unit_0_alu_0_n_14_9),.ZN(execution_unit_0_alu_0_n_57));
	INV_X1_LVT execution_unit_0alu_0i_15_0 (.A(execution_unit_0_alu_0_n_57),.ZN(execution_unit_0_alu_0_n_58));
	HA_X1_LVT execution_unit_0alu_0i_16_0 (.A(execution_unit_0_alu_0_n_52),.B(execution_unit_0_alu_0_n_53),.CO(execution_unit_0_alu_0_n_16_0),.S(execution_unit_0_alu_0_n_59));
	FA_X1_LVT execution_unit_0alu_0i_16_1 (.A(execution_unit_0_alu_0_n_55),.B(execution_unit_0_alu_0_n_54),.CI(execution_unit_0_alu_0_n_16_0),.CO(execution_unit_0_alu_0_n_16_1),.S(execution_unit_0_alu_0_n_60));
	OR2_X1_LVT execution_unit_0alu_0i_17_7 (.A1(execution_unit_0_alu_0_n_58),.A2(execution_unit_0_alu_0_n_60),.ZN(execution_unit_0_alu_0_n_17_5));
	HA_X1_LVT execution_unit_0alu_0i_16_2 (.A(execution_unit_0_alu_0_n_56),.B(execution_unit_0_alu_0_n_16_1),.CO(execution_unit_0_alu_0_n_16_2),.S(execution_unit_0_alu_0_n_61));
	INV_X1_LVT execution_unit_0alu_0i_17_8 (.A(execution_unit_0_alu_0_n_61),.ZN(execution_unit_0_alu_0_n_17_6));
	XNOR2_X1_LVT execution_unit_0alu_0i_17_10 (.A(execution_unit_0_alu_0_n_17_5),.B(execution_unit_0_alu_0_n_17_6),.ZN(execution_unit_0_alu_0_n_17_8));
	INV_X1_LVT execution_unit_0alu_0i_17_3 (.A(execution_unit_0_alu_0_n_51),.ZN(execution_unit_0_alu_0_n_17_2));
	NAND2_X1_LVT execution_unit_0alu_0i_17_2 (.A1(execution_unit_0_alu_0_n_58),.A2(execution_unit_0_alu_0_n_17_2),.ZN(execution_unit_0_alu_0_n_17_1));
	OR2_X1_LVT execution_unit_0alu_0i_17_5 (.A1(execution_unit_0_alu_0_n_59),.A2(execution_unit_0_alu_0_n_17_1),.ZN(execution_unit_0_alu_0_n_17_3));
	XNOR2_X1_LVT execution_unit_0alu_0i_17_6 (.A(execution_unit_0_alu_0_n_58),.B(execution_unit_0_alu_0_n_60),.ZN(execution_unit_0_alu_0_n_17_4));
	HA_X1_LVT execution_unit_0alu_0i_17_9 (.A(execution_unit_0_alu_0_n_17_3),.B(execution_unit_0_alu_0_n_17_4),.CO(execution_unit_0_alu_0_n_17_7),.S(execution_unit_0_alu_0_bcd_add0[3]));
	XNOR2_X1_LVT execution_unit_0alu_0i_17_11 (.A(execution_unit_0_alu_0_n_17_8),.B(execution_unit_0_alu_0_n_17_7),.ZN(execution_unit_0_alu_0_bcd_add0[4]));
	FA_X1_LVT execution_unit_0alu_0i_18_0 (.A(execution_unit_0_alu_0_n_0),.B(execution_unit_0_alu_0_bcd_add0[4]),.CI(execution_unit_0_alu_0_n_16),.CO(execution_unit_0_alu_0_n_18_0),.S(execution_unit_0_alu_0_n_62));
	FA_X1_LVT execution_unit_0alu_0i_18_1 (.A(execution_unit_0_alu_0_n_1),.B(execution_unit_0_alu_0_n_17),.CI(execution_unit_0_alu_0_n_18_0),.CO(execution_unit_0_alu_0_n_64),.S(execution_unit_0_alu_0_n_63));
	INV_X1_LVT execution_unit_0alu_0i_19_0 (.A(execution_unit_0_alu_0_n_64),.ZN(execution_unit_0_alu_0_n_19_0));
	FA_X1_LVT execution_unit_0alu_0i_19_3 (.A(execution_unit_0_alu_0_n_65),.B(execution_unit_0_alu_0_n_19_0),.CI(execution_unit_0_alu_0_n_63),.CO(execution_unit_0_alu_0_n_19_4),.S());
	FA_X1_LVT execution_unit_0alu_0i_19_4 (.A(execution_unit_0_alu_0_n_64),.B(execution_unit_0_alu_0_n_19_1),.CI(execution_unit_0_alu_0_n_19_4),.CO(execution_unit_0_alu_0_n_19_5),.S());
	FA_X1_LVT execution_unit_0alu_0i_19_5 (.A(execution_unit_0_alu_0_n_19_2),.B(execution_unit_0_alu_0_n_19_3),.CI(execution_unit_0_alu_0_n_19_5),.CO(execution_unit_0_alu_0_n_19_6),.S());
	HA_X1_LVT execution_unit_0alu_0i_19_6 (.A(execution_unit_0_alu_0_n_19_3),.B(execution_unit_0_alu_0_n_19_6),.CO(execution_unit_0_alu_0_n_19_7),.S());
	HA_X1_LVT execution_unit_0alu_0i_19_7 (.A(execution_unit_0_alu_0_n_19_3),.B(execution_unit_0_alu_0_n_19_7),.CO(execution_unit_0_alu_0_n_19_8),.S());
	XNOR2_X1_LVT execution_unit_0alu_0i_19_8 (.A(execution_unit_0_alu_0_n_19_3),.B(execution_unit_0_alu_0_n_19_8),.ZN(execution_unit_0_alu_0_n_19_9));
	INV_X1_LVT execution_unit_0alu_0i_19_9 (.A(execution_unit_0_alu_0_n_19_9),.ZN(execution_unit_0_alu_0_n_69));
	INV_X1_LVT execution_unit_0alu_0i_20_0 (.A(execution_unit_0_alu_0_n_69),.ZN(execution_unit_0_alu_0_n_70));
	HA_X1_LVT execution_unit_0alu_0i_21_0 (.A(execution_unit_0_alu_0_n_64),.B(execution_unit_0_alu_0_n_65),.CO(execution_unit_0_alu_0_n_21_0),.S(execution_unit_0_alu_0_n_71));
	FA_X1_LVT execution_unit_0alu_0i_21_1 (.A(execution_unit_0_alu_0_n_67),.B(execution_unit_0_alu_0_n_66),.CI(execution_unit_0_alu_0_n_21_0),.CO(execution_unit_0_alu_0_n_21_1),.S(execution_unit_0_alu_0_n_72));
	OR2_X1_LVT execution_unit_0alu_0i_22_7 (.A1(execution_unit_0_alu_0_n_70),.A2(execution_unit_0_alu_0_n_72),.ZN(execution_unit_0_alu_0_n_22_5));
	HA_X1_LVT execution_unit_0alu_0i_21_2 (.A(execution_unit_0_alu_0_n_68),.B(execution_unit_0_alu_0_n_21_1),.CO(execution_unit_0_alu_0_n_21_2),.S(execution_unit_0_alu_0_n_73));
	INV_X1_LVT execution_unit_0alu_0i_22_8 (.A(execution_unit_0_alu_0_n_73),.ZN(execution_unit_0_alu_0_n_22_6));
	XNOR2_X1_LVT execution_unit_0alu_0i_22_10 (.A(execution_unit_0_alu_0_n_22_5),.B(execution_unit_0_alu_0_n_22_6),.ZN(execution_unit_0_alu_0_n_22_8));
	INV_X1_LVT execution_unit_0alu_0i_22_3 (.A(execution_unit_0_alu_0_n_63),.ZN(execution_unit_0_alu_0_n_22_2));
	NAND2_X1_LVT execution_unit_0alu_0i_22_2 (.A1(execution_unit_0_alu_0_n_70),.A2(execution_unit_0_alu_0_n_22_2),.ZN(execution_unit_0_alu_0_n_22_1));
	OR2_X1_LVT execution_unit_0alu_0i_22_5 (.A1(execution_unit_0_alu_0_n_71),.A2(execution_unit_0_alu_0_n_22_1),.ZN(execution_unit_0_alu_0_n_22_3));
	XNOR2_X1_LVT execution_unit_0alu_0i_22_6 (.A(execution_unit_0_alu_0_n_70),.B(execution_unit_0_alu_0_n_72),.ZN(execution_unit_0_alu_0_n_22_4));
	HA_X1_LVT execution_unit_0alu_0i_22_9 (.A(execution_unit_0_alu_0_n_22_3),.B(execution_unit_0_alu_0_n_22_4),.CO(execution_unit_0_alu_0_n_22_7),.S(execution_unit_0_alu_0_bcd_add1[3]));
	XNOR2_X1_LVT execution_unit_0alu_0i_22_11 (.A(execution_unit_0_alu_0_n_22_8),.B(execution_unit_0_alu_0_n_22_7),.ZN(execution_unit_0_alu_0_bcd_add1[4]));
	FA_X1_LVT execution_unit_0alu_0i_23_0 (.A(execution_unit_0_alu_0_n_4),.B(execution_unit_0_alu_0_bcd_add1[4]),.CI(execution_unit_0_alu_0_X[0]),.CO(execution_unit_0_alu_0_n_23_0),.S(execution_unit_0_alu_0_n_74));
	FA_X1_LVT execution_unit_0alu_0i_23_1 (.A(execution_unit_0_alu_0_n_5),.B(execution_unit_0_alu_0_X[1]),.CI(execution_unit_0_alu_0_n_23_0),.CO(execution_unit_0_alu_0_n_76),.S(execution_unit_0_alu_0_n_75));
	HA_X1_LVT execution_unit_0alu_0i_23_2 (.A(execution_unit_0_alu_0_n_6),.B(execution_unit_0_alu_0_X[2]),.CO(execution_unit_0_alu_0_n_78),.S(execution_unit_0_alu_0_n_77));
	HA_X1_LVT execution_unit_0alu_0i_26_0 (.A(execution_unit_0_alu_0_n_76),.B(execution_unit_0_alu_0_n_77),.CO(execution_unit_0_alu_0_n_26_0),.S(execution_unit_0_alu_0_n_83));
	HA_X1_LVT execution_unit_0alu_0i_23_3 (.A(execution_unit_0_alu_0_n_7),.B(execution_unit_0_alu_0_X[3]),.CO(execution_unit_0_alu_0_n_80),.S(execution_unit_0_alu_0_n_79));
	INV_X1_LVT execution_unit_0alu_0i_24_2 (.A(execution_unit_0_alu_0_n_80),.ZN(execution_unit_0_alu_0_n_24_3));
	HA_X1_LVT execution_unit_0alu_0i_24_1 (.A(execution_unit_0_alu_0_n_79),.B(execution_unit_0_alu_0_n_78),.CO(execution_unit_0_alu_0_n_24_2),.S(execution_unit_0_alu_0_n_24_1));
	INV_X1_LVT execution_unit_0alu_0i_24_0 (.A(execution_unit_0_alu_0_n_76),.ZN(execution_unit_0_alu_0_n_24_0));
	FA_X1_LVT execution_unit_0alu_0i_24_3 (.A(execution_unit_0_alu_0_n_77),.B(execution_unit_0_alu_0_n_24_0),.CI(execution_unit_0_alu_0_n_75),.CO(execution_unit_0_alu_0_n_24_4),.S());
	FA_X1_LVT execution_unit_0alu_0i_24_4 (.A(execution_unit_0_alu_0_n_76),.B(execution_unit_0_alu_0_n_24_1),.CI(execution_unit_0_alu_0_n_24_4),.CO(execution_unit_0_alu_0_n_24_5),.S());
	FA_X1_LVT execution_unit_0alu_0i_24_5 (.A(execution_unit_0_alu_0_n_24_2),.B(execution_unit_0_alu_0_n_24_3),.CI(execution_unit_0_alu_0_n_24_5),.CO(execution_unit_0_alu_0_n_24_6),.S());
	HA_X1_LVT execution_unit_0alu_0i_24_6 (.A(execution_unit_0_alu_0_n_24_3),.B(execution_unit_0_alu_0_n_24_6),.CO(execution_unit_0_alu_0_n_24_7),.S());
	HA_X1_LVT execution_unit_0alu_0i_24_7 (.A(execution_unit_0_alu_0_n_24_3),.B(execution_unit_0_alu_0_n_24_7),.CO(execution_unit_0_alu_0_n_24_8),.S());
	XNOR2_X1_LVT execution_unit_0alu_0i_24_8 (.A(execution_unit_0_alu_0_n_24_3),.B(execution_unit_0_alu_0_n_24_8),.ZN(execution_unit_0_alu_0_n_24_9));
	INV_X1_LVT execution_unit_0alu_0i_24_9 (.A(execution_unit_0_alu_0_n_24_9),.ZN(execution_unit_0_alu_0_n_81));
	INV_X1_LVT execution_unit_0alu_0i_25_0 (.A(execution_unit_0_alu_0_n_81),.ZN(execution_unit_0_alu_0_n_82));
	INV_X1_LVT execution_unit_0alu_0i_27_3 (.A(execution_unit_0_alu_0_n_75),.ZN(execution_unit_0_alu_0_n_27_2));
	NAND2_X1_LVT execution_unit_0alu_0i_27_2 (.A1(execution_unit_0_alu_0_n_82),.A2(execution_unit_0_alu_0_n_27_2),.ZN(execution_unit_0_alu_0_n_27_1));
	OR2_X1_LVT execution_unit_0alu_0i_27_5 (.A1(execution_unit_0_alu_0_n_83),.A2(execution_unit_0_alu_0_n_27_1),.ZN(execution_unit_0_alu_0_n_27_3));
	FA_X1_LVT execution_unit_0alu_0i_26_1 (.A(execution_unit_0_alu_0_n_79),.B(execution_unit_0_alu_0_n_78),.CI(execution_unit_0_alu_0_n_26_0),.CO(execution_unit_0_alu_0_n_26_1),.S(execution_unit_0_alu_0_n_84));
	XNOR2_X1_LVT execution_unit_0alu_0i_27_6 (.A(execution_unit_0_alu_0_n_82),.B(execution_unit_0_alu_0_n_84),.ZN(execution_unit_0_alu_0_n_27_4));
	HA_X1_LVT execution_unit_0alu_0i_27_9 (.A(execution_unit_0_alu_0_n_27_3),.B(execution_unit_0_alu_0_n_27_4),.CO(execution_unit_0_alu_0_n_27_7),.S(execution_unit_0_alu_0_bcd_add2[3]));
	NOR2_X1_LVT execution_unit_0alu_0i_43_0 (.A1(inst_alu[7]),.A2(execution_unit_0_alu_0_n_104),.ZN(execution_unit_0_alu_0_n_105));
	OR4_X1_LVT execution_unit_0alu_0i_6_0 (.A1(inst_so[1]),.A2(inst_alu[10]),.A3(inst_alu[6]),.A4(inst_alu[5]),.ZN(execution_unit_0_alu_0_n_6_0));
	NOR3_X1_LVT execution_unit_0alu_0i_6_1 (.A1(execution_unit_0_alu_0_n_6_0),.A2(inst_alu[4]),.A3(inst_so[3]),.ZN(execution_unit_0_alu_0_alu_short_thro));
	NAND2_X1_LVT execution_unit_0alu_0i_7_143 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_X[3]),.ZN(execution_unit_0_alu_0_n_7_128));
	NAND2_X1_LVT execution_unit_0alu_0i_7_71 (.A1(inst_so[3]),.A2(execution_unit_0_n_117),.ZN(execution_unit_0_alu_0_n_7_64));
	NAND2_X1_LVT execution_unit_0alu_0i_7_144 (.A1(inst_so[1]),.A2(execution_unit_0_n_117),.ZN(execution_unit_0_alu_0_n_7_129));
	INV_X1_LVT execution_unit_0alu_0i_5_0 (.A(inst_bw),.ZN(execution_unit_0_alu_0_n_5_0));
	INV_X1_LVT execution_unit_0alu_0i_5_1 (.A(inst_so[0]),.ZN(execution_unit_0_alu_0_n_5_1));
	NAND3_X1_LVT execution_unit_0alu_0i_5_2 (.A1(execution_unit_0_alu_0_n_5_0),.A2(execution_unit_0_alu_0_n_5_1),.A3(execution_unit_0_n_109),.ZN(execution_unit_0_alu_0_n_5_2));
	NAND3_X1_LVT execution_unit_0alu_0i_5_3 (.A1(execution_unit_0_alu_0_n_5_1),.A2(inst_bw),.A3(execution_unit_0_n_117),.ZN(execution_unit_0_alu_0_n_5_3));
	NAND2_X1_LVT execution_unit_0alu_0i_5_4 (.A1(execution_unit_0_status[0]),.A2(inst_so[0]),.ZN(execution_unit_0_alu_0_n_5_4));
	NAND3_X1_LVT execution_unit_0alu_0i_5_5 (.A1(execution_unit_0_alu_0_n_5_2),.A2(execution_unit_0_alu_0_n_5_3),.A3(execution_unit_0_alu_0_n_5_4),.ZN(execution_unit_0_alu_0_n_20));
	NAND2_X1_LVT execution_unit_0alu_0i_7_145 (.A1(inst_alu[10]),.A2(execution_unit_0_alu_0_n_20),.ZN(execution_unit_0_alu_0_n_7_130));
	AND4_X1_LVT execution_unit_0alu_0i_7_146 (.A1(execution_unit_0_alu_0_n_7_128),.A2(execution_unit_0_alu_0_n_7_64),.A3(execution_unit_0_alu_0_n_7_129),.A4(execution_unit_0_alu_0_n_7_130),.ZN(execution_unit_0_alu_0_n_7_131));
	OAI21_X1_LVT execution_unit_0alu_0i_7_147 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_X[3]),.B2(execution_unit_0_alu_0_n_7),.ZN(execution_unit_0_alu_0_n_7_132));
	XOR2_X1_LVT execution_unit_0alu_0i_7_148 (.A(execution_unit_0_alu_0_X[3]),.B(execution_unit_0_alu_0_n_7),.Z(execution_unit_0_alu_0_n_7_133));
	NAND2_X1_LVT execution_unit_0alu_0i_7_149 (.A1(execution_unit_0_alu_0_n_7_133),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_134));
	NAND3_X1_LVT execution_unit_0alu_0i_7_150 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_X[3]),.A3(execution_unit_0_alu_0_n_7),.ZN(execution_unit_0_alu_0_n_7_135));
	NAND4_X1_LVT execution_unit_0alu_0i_7_151 (.A1(execution_unit_0_alu_0_n_7_131),.A2(execution_unit_0_alu_0_n_7_132),.A3(execution_unit_0_alu_0_n_7_134),.A4(execution_unit_0_alu_0_n_7_135),.ZN(execution_unit_0_alu_0_n_37));
	AOI222_X1_LVT execution_unit_0alu_0i_44_30 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[15]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add2[3]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_37),.ZN(execution_unit_0_alu_0_n_44_15));
	INV_X1_LVT execution_unit_0alu_0i_44_31 (.A(execution_unit_0_alu_0_n_44_15),.ZN(execution_unit_0_alu_out[15]));
	XNOR2_X1_LVT execution_unit_0alu_0i_27_4 (.A(execution_unit_0_alu_0_n_83),.B(execution_unit_0_alu_0_n_27_1),.ZN(execution_unit_0_alu_0_bcd_add2[2]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_134 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_X[2]),.ZN(execution_unit_0_alu_0_n_7_120));
	NAND2_X1_LVT execution_unit_0alu_0i_7_135 (.A1(inst_so[1]),.A2(execution_unit_0_n_118),.ZN(execution_unit_0_alu_0_n_7_121));
	NAND2_X1_LVT execution_unit_0alu_0i_7_136 (.A1(inst_alu[10]),.A2(execution_unit_0_n_109),.ZN(execution_unit_0_alu_0_n_7_122));
	AND4_X1_LVT execution_unit_0alu_0i_7_137 (.A1(execution_unit_0_alu_0_n_7_120),.A2(execution_unit_0_alu_0_n_7_64),.A3(execution_unit_0_alu_0_n_7_121),.A4(execution_unit_0_alu_0_n_7_122),.ZN(execution_unit_0_alu_0_n_7_123));
	OAI21_X1_LVT execution_unit_0alu_0i_7_138 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_X[2]),.B2(execution_unit_0_alu_0_n_6),.ZN(execution_unit_0_alu_0_n_7_124));
	XOR2_X1_LVT execution_unit_0alu_0i_7_139 (.A(execution_unit_0_alu_0_X[2]),.B(execution_unit_0_alu_0_n_6),.Z(execution_unit_0_alu_0_n_7_125));
	NAND2_X1_LVT execution_unit_0alu_0i_7_140 (.A1(execution_unit_0_alu_0_n_7_125),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_126));
	NAND3_X1_LVT execution_unit_0alu_0i_7_141 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_X[2]),.A3(execution_unit_0_alu_0_n_6),.ZN(execution_unit_0_alu_0_n_7_127));
	NAND4_X1_LVT execution_unit_0alu_0i_7_142 (.A1(execution_unit_0_alu_0_n_7_123),.A2(execution_unit_0_alu_0_n_7_124),.A3(execution_unit_0_alu_0_n_7_126),.A4(execution_unit_0_alu_0_n_7_127),.ZN(execution_unit_0_alu_0_n_36));
	AOI222_X1_LVT execution_unit_0alu_0i_44_28 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[14]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add2[2]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_36),.ZN(execution_unit_0_alu_0_n_44_14));
	INV_X1_LVT execution_unit_0alu_0i_44_29 (.A(execution_unit_0_alu_0_n_44_14),.ZN(execution_unit_0_alu_out[14]));
	XNOR2_X1_LVT execution_unit_0alu_0i_27_0 (.A(execution_unit_0_alu_0_n_82),.B(execution_unit_0_alu_0_n_75),.ZN(execution_unit_0_alu_0_n_27_0));
	INV_X1_LVT execution_unit_0alu_0i_27_1 (.A(execution_unit_0_alu_0_n_27_0),.ZN(execution_unit_0_alu_0_bcd_add2[1]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_125 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_X[1]),.ZN(execution_unit_0_alu_0_n_7_112));
	NAND2_X1_LVT execution_unit_0alu_0i_7_126 (.A1(inst_so[1]),.A2(execution_unit_0_n_119),.ZN(execution_unit_0_alu_0_n_7_113));
	NAND2_X1_LVT execution_unit_0alu_0i_7_127 (.A1(inst_alu[10]),.A2(execution_unit_0_n_110),.ZN(execution_unit_0_alu_0_n_7_114));
	AND4_X1_LVT execution_unit_0alu_0i_7_128 (.A1(execution_unit_0_alu_0_n_7_112),.A2(execution_unit_0_alu_0_n_7_64),.A3(execution_unit_0_alu_0_n_7_113),.A4(execution_unit_0_alu_0_n_7_114),.ZN(execution_unit_0_alu_0_n_7_115));
	OAI21_X1_LVT execution_unit_0alu_0i_7_129 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_X[1]),.B2(execution_unit_0_alu_0_n_5),.ZN(execution_unit_0_alu_0_n_7_116));
	XOR2_X1_LVT execution_unit_0alu_0i_7_130 (.A(execution_unit_0_alu_0_X[1]),.B(execution_unit_0_alu_0_n_5),.Z(execution_unit_0_alu_0_n_7_117));
	NAND2_X1_LVT execution_unit_0alu_0i_7_131 (.A1(execution_unit_0_alu_0_n_7_117),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_118));
	NAND3_X1_LVT execution_unit_0alu_0i_7_132 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_X[1]),.A3(execution_unit_0_alu_0_n_5),.ZN(execution_unit_0_alu_0_n_7_119));
	NAND4_X1_LVT execution_unit_0alu_0i_7_133 (.A1(execution_unit_0_alu_0_n_7_115),.A2(execution_unit_0_alu_0_n_7_116),.A3(execution_unit_0_alu_0_n_7_118),.A4(execution_unit_0_alu_0_n_7_119),.ZN(execution_unit_0_alu_0_n_35));
	AOI222_X1_LVT execution_unit_0alu_0i_44_26 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[13]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add2[1]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_35),.ZN(execution_unit_0_alu_0_n_44_13));
	INV_X1_LVT execution_unit_0alu_0i_44_27 (.A(execution_unit_0_alu_0_n_44_13),.ZN(execution_unit_0_alu_out[13]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_116 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_X[0]),.ZN(execution_unit_0_alu_0_n_7_104));
	NAND2_X1_LVT execution_unit_0alu_0i_7_117 (.A1(inst_so[1]),.A2(execution_unit_0_n_120),.ZN(execution_unit_0_alu_0_n_7_105));
	NAND2_X1_LVT execution_unit_0alu_0i_7_118 (.A1(inst_alu[10]),.A2(execution_unit_0_n_111),.ZN(execution_unit_0_alu_0_n_7_106));
	AND4_X1_LVT execution_unit_0alu_0i_7_119 (.A1(execution_unit_0_alu_0_n_7_104),.A2(execution_unit_0_alu_0_n_7_64),.A3(execution_unit_0_alu_0_n_7_105),.A4(execution_unit_0_alu_0_n_7_106),.ZN(execution_unit_0_alu_0_n_7_107));
	OAI21_X1_LVT execution_unit_0alu_0i_7_120 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_X[0]),.B2(execution_unit_0_alu_0_n_4),.ZN(execution_unit_0_alu_0_n_7_108));
	XOR2_X1_LVT execution_unit_0alu_0i_7_121 (.A(execution_unit_0_alu_0_X[0]),.B(execution_unit_0_alu_0_n_4),.Z(execution_unit_0_alu_0_n_7_109));
	NAND2_X1_LVT execution_unit_0alu_0i_7_122 (.A1(execution_unit_0_alu_0_n_7_109),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_110));
	NAND3_X1_LVT execution_unit_0alu_0i_7_123 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_X[0]),.A3(execution_unit_0_alu_0_n_4),.ZN(execution_unit_0_alu_0_n_7_111));
	NAND4_X1_LVT execution_unit_0alu_0i_7_124 (.A1(execution_unit_0_alu_0_n_7_107),.A2(execution_unit_0_alu_0_n_7_108),.A3(execution_unit_0_alu_0_n_7_110),.A4(execution_unit_0_alu_0_n_7_111),.ZN(execution_unit_0_alu_0_n_34));
	AOI222_X1_LVT execution_unit_0alu_0i_44_24 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[12]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_n_74),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_34),.ZN(execution_unit_0_alu_0_n_44_12));
	INV_X1_LVT execution_unit_0alu_0i_44_25 (.A(execution_unit_0_alu_0_n_44_12),.ZN(execution_unit_0_alu_out[12]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_107 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_19),.ZN(execution_unit_0_alu_0_n_7_96));
	NAND2_X1_LVT execution_unit_0alu_0i_7_108 (.A1(inst_so[1]),.A2(execution_unit_0_n_121),.ZN(execution_unit_0_alu_0_n_7_97));
	NAND2_X1_LVT execution_unit_0alu_0i_7_109 (.A1(inst_alu[10]),.A2(execution_unit_0_n_112),.ZN(execution_unit_0_alu_0_n_7_98));
	AND4_X1_LVT execution_unit_0alu_0i_7_110 (.A1(execution_unit_0_alu_0_n_7_96),.A2(execution_unit_0_alu_0_n_7_64),.A3(execution_unit_0_alu_0_n_7_97),.A4(execution_unit_0_alu_0_n_7_98),.ZN(execution_unit_0_alu_0_n_7_99));
	OAI21_X1_LVT execution_unit_0alu_0i_7_111 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_19),.B2(execution_unit_0_alu_0_n_3),.ZN(execution_unit_0_alu_0_n_7_100));
	XOR2_X1_LVT execution_unit_0alu_0i_7_112 (.A(execution_unit_0_alu_0_n_19),.B(execution_unit_0_alu_0_n_3),.Z(execution_unit_0_alu_0_n_7_101));
	NAND2_X1_LVT execution_unit_0alu_0i_7_113 (.A1(execution_unit_0_alu_0_n_7_101),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_102));
	NAND3_X1_LVT execution_unit_0alu_0i_7_114 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_19),.A3(execution_unit_0_alu_0_n_3),.ZN(execution_unit_0_alu_0_n_7_103));
	NAND4_X1_LVT execution_unit_0alu_0i_7_115 (.A1(execution_unit_0_alu_0_n_7_99),.A2(execution_unit_0_alu_0_n_7_100),.A3(execution_unit_0_alu_0_n_7_102),.A4(execution_unit_0_alu_0_n_7_103),.ZN(execution_unit_0_alu_0_n_33));
	AOI222_X1_LVT execution_unit_0alu_0i_44_22 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[11]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add1[3]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_33),.ZN(execution_unit_0_alu_0_n_44_11));
	INV_X1_LVT execution_unit_0alu_0i_44_23 (.A(execution_unit_0_alu_0_n_44_11),.ZN(execution_unit_0_alu_out[11]));
	XNOR2_X1_LVT execution_unit_0alu_0i_22_4 (.A(execution_unit_0_alu_0_n_71),.B(execution_unit_0_alu_0_n_22_1),.ZN(execution_unit_0_alu_0_bcd_add1[2]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_98 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_18),.ZN(execution_unit_0_alu_0_n_7_88));
	NAND2_X1_LVT execution_unit_0alu_0i_7_99 (.A1(inst_so[1]),.A2(execution_unit_0_n_122),.ZN(execution_unit_0_alu_0_n_7_89));
	NAND2_X1_LVT execution_unit_0alu_0i_7_100 (.A1(inst_alu[10]),.A2(execution_unit_0_n_113),.ZN(execution_unit_0_alu_0_n_7_90));
	AND4_X1_LVT execution_unit_0alu_0i_7_101 (.A1(execution_unit_0_alu_0_n_7_88),.A2(execution_unit_0_alu_0_n_7_64),.A3(execution_unit_0_alu_0_n_7_89),.A4(execution_unit_0_alu_0_n_7_90),.ZN(execution_unit_0_alu_0_n_7_91));
	OAI21_X1_LVT execution_unit_0alu_0i_7_102 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_18),.B2(execution_unit_0_alu_0_n_2),.ZN(execution_unit_0_alu_0_n_7_92));
	XOR2_X1_LVT execution_unit_0alu_0i_7_103 (.A(execution_unit_0_alu_0_n_18),.B(execution_unit_0_alu_0_n_2),.Z(execution_unit_0_alu_0_n_7_93));
	NAND2_X1_LVT execution_unit_0alu_0i_7_104 (.A1(execution_unit_0_alu_0_n_7_93),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_94));
	NAND3_X1_LVT execution_unit_0alu_0i_7_105 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_18),.A3(execution_unit_0_alu_0_n_2),.ZN(execution_unit_0_alu_0_n_7_95));
	NAND4_X1_LVT execution_unit_0alu_0i_7_106 (.A1(execution_unit_0_alu_0_n_7_91),.A2(execution_unit_0_alu_0_n_7_92),.A3(execution_unit_0_alu_0_n_7_94),.A4(execution_unit_0_alu_0_n_7_95),.ZN(execution_unit_0_alu_0_n_32));
	AOI222_X1_LVT execution_unit_0alu_0i_44_20 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[10]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add1[2]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_32),.ZN(execution_unit_0_alu_0_n_44_10));
	INV_X1_LVT execution_unit_0alu_0i_44_21 (.A(execution_unit_0_alu_0_n_44_10),.ZN(execution_unit_0_alu_out[10]));
	XNOR2_X1_LVT execution_unit_0alu_0i_22_0 (.A(execution_unit_0_alu_0_n_70),.B(execution_unit_0_alu_0_n_63),.ZN(execution_unit_0_alu_0_n_22_0));
	INV_X1_LVT execution_unit_0alu_0i_22_1 (.A(execution_unit_0_alu_0_n_22_0),.ZN(execution_unit_0_alu_0_bcd_add1[1]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_89 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_17),.ZN(execution_unit_0_alu_0_n_7_80));
	NAND2_X1_LVT execution_unit_0alu_0i_7_90 (.A1(inst_so[1]),.A2(execution_unit_0_n_123),.ZN(execution_unit_0_alu_0_n_7_81));
	NAND2_X1_LVT execution_unit_0alu_0i_7_91 (.A1(inst_alu[10]),.A2(execution_unit_0_n_114),.ZN(execution_unit_0_alu_0_n_7_82));
	AND4_X1_LVT execution_unit_0alu_0i_7_92 (.A1(execution_unit_0_alu_0_n_7_80),.A2(execution_unit_0_alu_0_n_7_64),.A3(execution_unit_0_alu_0_n_7_81),.A4(execution_unit_0_alu_0_n_7_82),.ZN(execution_unit_0_alu_0_n_7_83));
	OAI21_X1_LVT execution_unit_0alu_0i_7_93 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_17),.B2(execution_unit_0_alu_0_n_1),.ZN(execution_unit_0_alu_0_n_7_84));
	XOR2_X1_LVT execution_unit_0alu_0i_7_94 (.A(execution_unit_0_alu_0_n_17),.B(execution_unit_0_alu_0_n_1),.Z(execution_unit_0_alu_0_n_7_85));
	NAND2_X1_LVT execution_unit_0alu_0i_7_95 (.A1(execution_unit_0_alu_0_n_7_85),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_86));
	NAND3_X1_LVT execution_unit_0alu_0i_7_96 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_17),.A3(execution_unit_0_alu_0_n_1),.ZN(execution_unit_0_alu_0_n_7_87));
	NAND4_X1_LVT execution_unit_0alu_0i_7_97 (.A1(execution_unit_0_alu_0_n_7_83),.A2(execution_unit_0_alu_0_n_7_84),.A3(execution_unit_0_alu_0_n_7_86),.A4(execution_unit_0_alu_0_n_7_87),.ZN(execution_unit_0_alu_0_n_31));
	AOI222_X1_LVT execution_unit_0alu_0i_44_18 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[9]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add1[1]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_31),.ZN(execution_unit_0_alu_0_n_44_9));
	INV_X1_LVT execution_unit_0alu_0i_44_19 (.A(execution_unit_0_alu_0_n_44_9),.ZN(execution_unit_0_alu_out[9]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_80 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_16),.ZN(execution_unit_0_alu_0_n_7_72));
	NAND2_X1_LVT execution_unit_0alu_0i_7_81 (.A1(execution_unit_0_n_124),.A2(inst_so[1]),.ZN(execution_unit_0_alu_0_n_7_73));
	NAND2_X1_LVT execution_unit_0alu_0i_7_82 (.A1(inst_alu[10]),.A2(execution_unit_0_n_115),.ZN(execution_unit_0_alu_0_n_7_74));
	AND4_X1_LVT execution_unit_0alu_0i_7_83 (.A1(execution_unit_0_alu_0_n_7_72),.A2(execution_unit_0_alu_0_n_7_64),.A3(execution_unit_0_alu_0_n_7_73),.A4(execution_unit_0_alu_0_n_7_74),.ZN(execution_unit_0_alu_0_n_7_75));
	OAI21_X1_LVT execution_unit_0alu_0i_7_84 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_16),.B2(execution_unit_0_alu_0_n_0),.ZN(execution_unit_0_alu_0_n_7_76));
	XOR2_X1_LVT execution_unit_0alu_0i_7_85 (.A(execution_unit_0_alu_0_n_16),.B(execution_unit_0_alu_0_n_0),.Z(execution_unit_0_alu_0_n_7_77));
	NAND2_X1_LVT execution_unit_0alu_0i_7_86 (.A1(execution_unit_0_alu_0_n_7_77),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_78));
	NAND3_X1_LVT execution_unit_0alu_0i_7_87 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_16),.A3(execution_unit_0_alu_0_n_0),.ZN(execution_unit_0_alu_0_n_7_79));
	NAND4_X1_LVT execution_unit_0alu_0i_7_88 (.A1(execution_unit_0_alu_0_n_7_75),.A2(execution_unit_0_alu_0_n_7_76),.A3(execution_unit_0_alu_0_n_7_78),.A4(execution_unit_0_alu_0_n_7_79),.ZN(execution_unit_0_alu_0_n_30));
	AOI222_X1_LVT execution_unit_0alu_0i_44_16 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[8]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_n_62),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_30),.ZN(execution_unit_0_alu_0_n_44_8));
	INV_X1_LVT execution_unit_0alu_0i_44_17 (.A(execution_unit_0_alu_0_n_44_8),.ZN(execution_unit_0_alu_out[8]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_70 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_15),.ZN(execution_unit_0_alu_0_n_7_63));
	NAND2_X1_LVT execution_unit_0alu_0i_7_72 (.A1(inst_so[1]),.A2(execution_unit_0_n_109),.ZN(execution_unit_0_alu_0_n_7_65));
	AOI22_X1_LVT execution_unit_0alu_0i_5_6 (.A1(execution_unit_0_alu_0_n_20),.A2(inst_bw),.B1(execution_unit_0_alu_0_n_5_0),.B2(execution_unit_0_n_116),.ZN(execution_unit_0_alu_0_n_5_5));
	INV_X1_LVT execution_unit_0alu_0i_5_7 (.A(execution_unit_0_alu_0_n_5_5),.ZN(execution_unit_0_alu_0_n_21));
	NAND2_X1_LVT execution_unit_0alu_0i_7_73 (.A1(inst_alu[10]),.A2(execution_unit_0_alu_0_n_21),.ZN(execution_unit_0_alu_0_n_7_66));
	AND4_X1_LVT execution_unit_0alu_0i_7_74 (.A1(execution_unit_0_alu_0_n_7_63),.A2(execution_unit_0_alu_0_n_7_64),.A3(execution_unit_0_alu_0_n_7_65),.A4(execution_unit_0_alu_0_n_7_66),.ZN(execution_unit_0_alu_0_n_7_67));
	OAI21_X1_LVT execution_unit_0alu_0i_7_75 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_15),.B2(execution_unit_0_n_86),.ZN(execution_unit_0_alu_0_n_7_68));
	XOR2_X1_LVT execution_unit_0alu_0i_7_76 (.A(execution_unit_0_alu_0_n_15),.B(execution_unit_0_n_86),.Z(execution_unit_0_alu_0_n_7_69));
	NAND2_X1_LVT execution_unit_0alu_0i_7_77 (.A1(execution_unit_0_alu_0_n_7_69),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_70));
	NAND3_X1_LVT execution_unit_0alu_0i_7_78 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_15),.A3(execution_unit_0_n_86),.ZN(execution_unit_0_alu_0_n_7_71));
	NAND4_X1_LVT execution_unit_0alu_0i_7_79 (.A1(execution_unit_0_alu_0_n_7_67),.A2(execution_unit_0_alu_0_n_7_68),.A3(execution_unit_0_alu_0_n_7_70),.A4(execution_unit_0_alu_0_n_7_71),.ZN(execution_unit_0_alu_0_n_29));
	AOI222_X1_LVT execution_unit_0alu_0i_44_14 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[7]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add0[3]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_29),.ZN(execution_unit_0_alu_0_n_44_7));
	INV_X1_LVT execution_unit_0alu_0i_44_15 (.A(execution_unit_0_alu_0_n_44_7),.ZN(execution_unit_0_alu_out[7]));
	XNOR2_X1_LVT execution_unit_0alu_0i_17_4 (.A(execution_unit_0_alu_0_n_59),.B(execution_unit_0_alu_0_n_17_1),.ZN(execution_unit_0_alu_0_bcd_add0[2]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_60 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_14),.ZN(execution_unit_0_alu_0_n_7_54));
	NAND2_X1_LVT execution_unit_0alu_0i_7_61 (.A1(inst_so[3]),.A2(execution_unit_0_n_118),.ZN(execution_unit_0_alu_0_n_7_55));
	NAND2_X1_LVT execution_unit_0alu_0i_7_62 (.A1(inst_so[1]),.A2(execution_unit_0_n_110),.ZN(execution_unit_0_alu_0_n_7_56));
	NAND2_X1_LVT execution_unit_0alu_0i_7_63 (.A1(inst_alu[10]),.A2(execution_unit_0_n_117),.ZN(execution_unit_0_alu_0_n_7_57));
	AND4_X1_LVT execution_unit_0alu_0i_7_64 (.A1(execution_unit_0_alu_0_n_7_54),.A2(execution_unit_0_alu_0_n_7_55),.A3(execution_unit_0_alu_0_n_7_56),.A4(execution_unit_0_alu_0_n_7_57),.ZN(execution_unit_0_alu_0_n_7_58));
	OAI21_X1_LVT execution_unit_0alu_0i_7_65 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_14),.B2(execution_unit_0_n_87),.ZN(execution_unit_0_alu_0_n_7_59));
	XOR2_X1_LVT execution_unit_0alu_0i_7_66 (.A(execution_unit_0_alu_0_n_14),.B(execution_unit_0_n_87),.Z(execution_unit_0_alu_0_n_7_60));
	NAND2_X1_LVT execution_unit_0alu_0i_7_67 (.A1(execution_unit_0_alu_0_n_7_60),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_61));
	NAND3_X1_LVT execution_unit_0alu_0i_7_68 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_14),.A3(execution_unit_0_n_87),.ZN(execution_unit_0_alu_0_n_7_62));
	NAND4_X1_LVT execution_unit_0alu_0i_7_69 (.A1(execution_unit_0_alu_0_n_7_58),.A2(execution_unit_0_alu_0_n_7_59),.A3(execution_unit_0_alu_0_n_7_61),.A4(execution_unit_0_alu_0_n_7_62),.ZN(execution_unit_0_alu_0_n_28));
	AOI222_X1_LVT execution_unit_0alu_0i_44_12 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[6]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add0[2]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_28),.ZN(execution_unit_0_alu_0_n_44_6));
	INV_X1_LVT execution_unit_0alu_0i_44_13 (.A(execution_unit_0_alu_0_n_44_6),.ZN(execution_unit_0_alu_out[6]));
	XNOR2_X1_LVT execution_unit_0alu_0i_17_0 (.A(execution_unit_0_alu_0_n_58),.B(execution_unit_0_alu_0_n_51),.ZN(execution_unit_0_alu_0_n_17_0));
	INV_X1_LVT execution_unit_0alu_0i_17_1 (.A(execution_unit_0_alu_0_n_17_0),.ZN(execution_unit_0_alu_0_bcd_add0[1]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_50 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_13),.ZN(execution_unit_0_alu_0_n_7_45));
	NAND2_X1_LVT execution_unit_0alu_0i_7_51 (.A1(inst_so[3]),.A2(execution_unit_0_n_119),.ZN(execution_unit_0_alu_0_n_7_46));
	NAND2_X1_LVT execution_unit_0alu_0i_7_52 (.A1(inst_so[1]),.A2(execution_unit_0_n_111),.ZN(execution_unit_0_alu_0_n_7_47));
	NAND2_X1_LVT execution_unit_0alu_0i_7_53 (.A1(inst_alu[10]),.A2(execution_unit_0_n_118),.ZN(execution_unit_0_alu_0_n_7_48));
	AND4_X1_LVT execution_unit_0alu_0i_7_54 (.A1(execution_unit_0_alu_0_n_7_45),.A2(execution_unit_0_alu_0_n_7_46),.A3(execution_unit_0_alu_0_n_7_47),.A4(execution_unit_0_alu_0_n_7_48),.ZN(execution_unit_0_alu_0_n_7_49));
	OAI21_X1_LVT execution_unit_0alu_0i_7_55 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_13),.B2(execution_unit_0_n_88),.ZN(execution_unit_0_alu_0_n_7_50));
	XOR2_X1_LVT execution_unit_0alu_0i_7_56 (.A(execution_unit_0_alu_0_n_13),.B(execution_unit_0_n_88),.Z(execution_unit_0_alu_0_n_7_51));
	NAND2_X1_LVT execution_unit_0alu_0i_7_57 (.A1(execution_unit_0_alu_0_n_7_51),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_52));
	NAND3_X1_LVT execution_unit_0alu_0i_7_58 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_13),.A3(execution_unit_0_n_88),.ZN(execution_unit_0_alu_0_n_7_53));
	NAND4_X1_LVT execution_unit_0alu_0i_7_59 (.A1(execution_unit_0_alu_0_n_7_49),.A2(execution_unit_0_alu_0_n_7_50),.A3(execution_unit_0_alu_0_n_7_52),.A4(execution_unit_0_alu_0_n_7_53),.ZN(execution_unit_0_alu_0_n_27));
	AOI222_X1_LVT execution_unit_0alu_0i_44_10 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[5]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add0[1]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_27),.ZN(execution_unit_0_alu_0_n_44_5));
	INV_X1_LVT execution_unit_0alu_0i_44_11 (.A(execution_unit_0_alu_0_n_44_5),.ZN(execution_unit_0_alu_out[5]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_40 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_12),.ZN(execution_unit_0_alu_0_n_7_36));
	NAND2_X1_LVT execution_unit_0alu_0i_7_41 (.A1(inst_so[3]),.A2(execution_unit_0_n_120),.ZN(execution_unit_0_alu_0_n_7_37));
	NAND2_X1_LVT execution_unit_0alu_0i_7_42 (.A1(inst_so[1]),.A2(execution_unit_0_n_112),.ZN(execution_unit_0_alu_0_n_7_38));
	NAND2_X1_LVT execution_unit_0alu_0i_7_43 (.A1(inst_alu[10]),.A2(execution_unit_0_n_119),.ZN(execution_unit_0_alu_0_n_7_39));
	AND4_X1_LVT execution_unit_0alu_0i_7_44 (.A1(execution_unit_0_alu_0_n_7_36),.A2(execution_unit_0_alu_0_n_7_37),.A3(execution_unit_0_alu_0_n_7_38),.A4(execution_unit_0_alu_0_n_7_39),.ZN(execution_unit_0_alu_0_n_7_40));
	OAI21_X1_LVT execution_unit_0alu_0i_7_45 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_12),.B2(execution_unit_0_n_89),.ZN(execution_unit_0_alu_0_n_7_41));
	XOR2_X1_LVT execution_unit_0alu_0i_7_46 (.A(execution_unit_0_alu_0_n_12),.B(execution_unit_0_n_89),.Z(execution_unit_0_alu_0_n_7_42));
	NAND2_X1_LVT execution_unit_0alu_0i_7_47 (.A1(execution_unit_0_alu_0_n_7_42),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_43));
	NAND3_X1_LVT execution_unit_0alu_0i_7_48 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_12),.A3(execution_unit_0_n_89),.ZN(execution_unit_0_alu_0_n_7_44));
	NAND4_X1_LVT execution_unit_0alu_0i_7_49 (.A1(execution_unit_0_alu_0_n_7_40),.A2(execution_unit_0_alu_0_n_7_41),.A3(execution_unit_0_alu_0_n_7_43),.A4(execution_unit_0_alu_0_n_7_44),.ZN(execution_unit_0_alu_0_n_26));
	AOI222_X1_LVT execution_unit_0alu_0i_44_8 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[4]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_n_50),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_26),.ZN(execution_unit_0_alu_0_n_44_4));
	INV_X1_LVT execution_unit_0alu_0i_44_9 (.A(execution_unit_0_alu_0_n_44_4),.ZN(execution_unit_0_alu_out[4]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_30 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_11),.ZN(execution_unit_0_alu_0_n_7_27));
	NAND2_X1_LVT execution_unit_0alu_0i_7_31 (.A1(inst_so[3]),.A2(execution_unit_0_n_121),.ZN(execution_unit_0_alu_0_n_7_28));
	NAND2_X1_LVT execution_unit_0alu_0i_7_32 (.A1(inst_so[1]),.A2(execution_unit_0_n_113),.ZN(execution_unit_0_alu_0_n_7_29));
	NAND2_X1_LVT execution_unit_0alu_0i_7_33 (.A1(inst_alu[10]),.A2(execution_unit_0_n_120),.ZN(execution_unit_0_alu_0_n_7_30));
	AND4_X1_LVT execution_unit_0alu_0i_7_34 (.A1(execution_unit_0_alu_0_n_7_27),.A2(execution_unit_0_alu_0_n_7_28),.A3(execution_unit_0_alu_0_n_7_29),.A4(execution_unit_0_alu_0_n_7_30),.ZN(execution_unit_0_alu_0_n_7_31));
	OAI21_X1_LVT execution_unit_0alu_0i_7_35 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_11),.B2(execution_unit_0_n_90),.ZN(execution_unit_0_alu_0_n_7_32));
	XOR2_X1_LVT execution_unit_0alu_0i_7_36 (.A(execution_unit_0_alu_0_n_11),.B(execution_unit_0_n_90),.Z(execution_unit_0_alu_0_n_7_33));
	NAND2_X1_LVT execution_unit_0alu_0i_7_37 (.A1(execution_unit_0_alu_0_n_7_33),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_34));
	NAND3_X1_LVT execution_unit_0alu_0i_7_38 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_11),.A3(execution_unit_0_n_90),.ZN(execution_unit_0_alu_0_n_7_35));
	NAND4_X1_LVT execution_unit_0alu_0i_7_39 (.A1(execution_unit_0_alu_0_n_7_31),.A2(execution_unit_0_alu_0_n_7_32),.A3(execution_unit_0_alu_0_n_7_34),.A4(execution_unit_0_alu_0_n_7_35),.ZN(execution_unit_0_alu_0_n_25));
	AOI222_X1_LVT execution_unit_0alu_0i_44_6 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[3]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add[3]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_25),.ZN(execution_unit_0_alu_0_n_44_3));
	INV_X1_LVT execution_unit_0alu_0i_44_7 (.A(execution_unit_0_alu_0_n_44_3),.ZN(execution_unit_0_alu_out[3]));
	XNOR2_X1_LVT execution_unit_0alu_0i_12_4 (.A(execution_unit_0_alu_0_n_47),.B(execution_unit_0_alu_0_n_12_1),.ZN(execution_unit_0_alu_0_bcd_add[2]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_20 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_10),.ZN(execution_unit_0_alu_0_n_7_18));
	NAND2_X1_LVT execution_unit_0alu_0i_7_21 (.A1(inst_so[3]),.A2(execution_unit_0_n_122),.ZN(execution_unit_0_alu_0_n_7_19));
	NAND2_X1_LVT execution_unit_0alu_0i_7_22 (.A1(inst_so[1]),.A2(execution_unit_0_n_114),.ZN(execution_unit_0_alu_0_n_7_20));
	NAND2_X1_LVT execution_unit_0alu_0i_7_23 (.A1(inst_alu[10]),.A2(execution_unit_0_n_121),.ZN(execution_unit_0_alu_0_n_7_21));
	AND4_X1_LVT execution_unit_0alu_0i_7_24 (.A1(execution_unit_0_alu_0_n_7_18),.A2(execution_unit_0_alu_0_n_7_19),.A3(execution_unit_0_alu_0_n_7_20),.A4(execution_unit_0_alu_0_n_7_21),.ZN(execution_unit_0_alu_0_n_7_22));
	OAI21_X1_LVT execution_unit_0alu_0i_7_25 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_10),.B2(execution_unit_0_n_91),.ZN(execution_unit_0_alu_0_n_7_23));
	XOR2_X1_LVT execution_unit_0alu_0i_7_26 (.A(execution_unit_0_alu_0_n_10),.B(execution_unit_0_n_91),.Z(execution_unit_0_alu_0_n_7_24));
	NAND2_X1_LVT execution_unit_0alu_0i_7_27 (.A1(execution_unit_0_alu_0_n_7_24),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_25));
	NAND3_X1_LVT execution_unit_0alu_0i_7_28 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_10),.A3(execution_unit_0_n_91),.ZN(execution_unit_0_alu_0_n_7_26));
	NAND4_X1_LVT execution_unit_0alu_0i_7_29 (.A1(execution_unit_0_alu_0_n_7_22),.A2(execution_unit_0_alu_0_n_7_23),.A3(execution_unit_0_alu_0_n_7_25),.A4(execution_unit_0_alu_0_n_7_26),.ZN(execution_unit_0_alu_0_n_24));
	AOI222_X1_LVT execution_unit_0alu_0i_44_4 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[2]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add[2]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_24),.ZN(execution_unit_0_alu_0_n_44_2));
	INV_X1_LVT execution_unit_0alu_0i_44_5 (.A(execution_unit_0_alu_0_n_44_2),.ZN(execution_unit_0_alu_out[2]));
	XNOR2_X1_LVT execution_unit_0alu_0i_12_0 (.A(execution_unit_0_alu_0_n_46),.B(execution_unit_0_alu_0_n_39),.ZN(execution_unit_0_alu_0_n_12_0));
	INV_X1_LVT execution_unit_0alu_0i_12_1 (.A(execution_unit_0_alu_0_n_12_0),.ZN(execution_unit_0_alu_0_bcd_add[1]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_10 (.A1(execution_unit_0_alu_0_alu_short_thro),.A2(execution_unit_0_alu_0_n_9),.ZN(execution_unit_0_alu_0_n_7_9));
	NAND2_X1_LVT execution_unit_0alu_0i_7_11 (.A1(inst_so[3]),.A2(execution_unit_0_n_123),.ZN(execution_unit_0_alu_0_n_7_10));
	NAND2_X1_LVT execution_unit_0alu_0i_7_12 (.A1(inst_so[1]),.A2(execution_unit_0_n_115),.ZN(execution_unit_0_alu_0_n_7_11));
	NAND2_X1_LVT execution_unit_0alu_0i_7_13 (.A1(inst_alu[10]),.A2(execution_unit_0_n_122),.ZN(execution_unit_0_alu_0_n_7_12));
	AND4_X1_LVT execution_unit_0alu_0i_7_14 (.A1(execution_unit_0_alu_0_n_7_9),.A2(execution_unit_0_alu_0_n_7_10),.A3(execution_unit_0_alu_0_n_7_11),.A4(execution_unit_0_alu_0_n_7_12),.ZN(execution_unit_0_alu_0_n_7_13));
	OAI21_X1_LVT execution_unit_0alu_0i_7_15 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_9),.B2(execution_unit_0_n_92),.ZN(execution_unit_0_alu_0_n_7_14));
	XOR2_X1_LVT execution_unit_0alu_0i_7_16 (.A(execution_unit_0_alu_0_n_9),.B(execution_unit_0_n_92),.Z(execution_unit_0_alu_0_n_7_15));
	NAND2_X1_LVT execution_unit_0alu_0i_7_17 (.A1(execution_unit_0_alu_0_n_7_15),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_16));
	NAND3_X1_LVT execution_unit_0alu_0i_7_18 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_9),.A3(execution_unit_0_n_92),.ZN(execution_unit_0_alu_0_n_7_17));
	NAND4_X1_LVT execution_unit_0alu_0i_7_19 (.A1(execution_unit_0_alu_0_n_7_13),.A2(execution_unit_0_alu_0_n_7_14),.A3(execution_unit_0_alu_0_n_7_16),.A4(execution_unit_0_alu_0_n_7_17),.ZN(execution_unit_0_alu_0_n_23));
	AOI222_X1_LVT execution_unit_0alu_0i_44_2 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[1]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add[1]),.C1(execution_unit_0_alu_0_n_105),.C2(execution_unit_0_alu_0_n_23),.ZN(execution_unit_0_alu_0_n_44_1));
	INV_X1_LVT execution_unit_0alu_0i_44_3 (.A(execution_unit_0_alu_0_n_44_1),.ZN(execution_unit_0_alu_out[1]));
	NAND2_X1_LVT execution_unit_0alu_0i_7_0 (.A1(execution_unit_0_alu_0_n_8),.A2(execution_unit_0_alu_0_alu_short_thro),.ZN(execution_unit_0_alu_0_n_7_0));
	NAND2_X1_LVT execution_unit_0alu_0i_7_1 (.A1(inst_so[3]),.A2(execution_unit_0_n_124),.ZN(execution_unit_0_alu_0_n_7_1));
	NAND2_X1_LVT execution_unit_0alu_0i_7_2 (.A1(inst_so[1]),.A2(execution_unit_0_n_116),.ZN(execution_unit_0_alu_0_n_7_2));
	NAND2_X1_LVT execution_unit_0alu_0i_7_3 (.A1(inst_alu[10]),.A2(execution_unit_0_n_123),.ZN(execution_unit_0_alu_0_n_7_3));
	AND4_X1_LVT execution_unit_0alu_0i_7_4 (.A1(execution_unit_0_alu_0_n_7_0),.A2(execution_unit_0_alu_0_n_7_1),.A3(execution_unit_0_alu_0_n_7_2),.A4(execution_unit_0_alu_0_n_7_3),.ZN(execution_unit_0_alu_0_n_7_4));
	OAI21_X1_LVT execution_unit_0alu_0i_7_5 (.A(inst_alu[5]),.B1(execution_unit_0_alu_0_n_8),.B2(execution_unit_0_n_93),.ZN(execution_unit_0_alu_0_n_7_5));
	XOR2_X1_LVT execution_unit_0alu_0i_7_6 (.A(execution_unit_0_alu_0_n_8),.B(execution_unit_0_n_93),.Z(execution_unit_0_alu_0_n_7_6));
	NAND2_X1_LVT execution_unit_0alu_0i_7_7 (.A1(execution_unit_0_alu_0_n_7_6),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_7_7));
	NAND3_X1_LVT execution_unit_0alu_0i_7_8 (.A1(inst_alu[4]),.A2(execution_unit_0_alu_0_n_8),.A3(execution_unit_0_n_93),.ZN(execution_unit_0_alu_0_n_7_8));
	NAND4_X1_LVT execution_unit_0alu_0i_7_9 (.A1(execution_unit_0_alu_0_n_7_4),.A2(execution_unit_0_alu_0_n_7_5),.A3(execution_unit_0_alu_0_n_7_7),.A4(execution_unit_0_alu_0_n_7_8),.ZN(execution_unit_0_alu_0_n_22));
	AOI222_X1_LVT execution_unit_0alu_0i_44_0 (.A1(execution_unit_0_alu_0_alu_add_inc[0]),.A2(execution_unit_0_alu_0_n_104),.B1(execution_unit_0_alu_0_n_38),.B2(execution_unit_0_alu_0_n_106),.C1(execution_unit_0_alu_0_n_22),.C2(execution_unit_0_alu_0_n_105),.ZN(execution_unit_0_alu_0_n_44_0));
	INV_X1_LVT execution_unit_0alu_0i_44_1 (.A(execution_unit_0_alu_0_n_44_0),.ZN(execution_unit_0_alu_out[0]));
	NOR2_X1_LVT execution_unit_0alu_0i_51_1 (.A1(inst_alu[8]),.A2(inst_alu[10]),.ZN(execution_unit_0_alu_0_n_51_1));
	NAND2_X1_LVT execution_unit_0alu_0i_51_2 (.A1(execution_unit_0_alu_0_n_51_1),.A2(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_51_2));
	INV_X1_LVT execution_unit_0alu_0i_51_8 (.A(inst_bw),.ZN(execution_unit_0_alu_0_n_51_8));
	AND2_X1_LVT execution_unit_0alu_0i_45_0 (.A1(execution_unit_0_alu_0_X[3]),.A2(execution_unit_0_alu_0_n_7),.ZN(execution_unit_0_alu_0_n_108));
	AND2_X1_LVT execution_unit_0alu_0i_47_0 (.A1(execution_unit_0_alu_0_n_15),.A2(execution_unit_0_n_86),.ZN(execution_unit_0_alu_0_n_110));
	AOI22_X1_LVT execution_unit_0alu_0i_51_24 (.A1(execution_unit_0_alu_0_n_51_8),.A2(execution_unit_0_alu_0_n_108),.B1(inst_bw),.B2(execution_unit_0_alu_0_n_110),.ZN(execution_unit_0_alu_0_n_51_21));
	INV_X1_LVT execution_unit_0alu_0i_51_6 (.A(inst_alu[6]),.ZN(execution_unit_0_alu_0_n_51_6));
	NAND2_X1_LVT execution_unit_0alu_0i_51_7 (.A1(execution_unit_0_alu_0_n_51_1),.A2(execution_unit_0_alu_0_n_51_6),.ZN(execution_unit_0_alu_0_n_51_7));
	INV_X1_LVT execution_unit_0alu_0i_46_0 (.A(execution_unit_0_alu_out[15]),.ZN(execution_unit_0_alu_0_n_46_0));
	NOR3_X1_LVT execution_unit_0alu_0i_46_1 (.A1(execution_unit_0_alu_0_n_46_0),.A2(execution_unit_0_alu_0_X[3]),.A3(execution_unit_0_alu_0_n_7),.ZN(execution_unit_0_alu_0_n_46_1));
	AOI21_X1_LVT execution_unit_0alu_0i_46_2 (.A(execution_unit_0_alu_0_n_46_1),.B1(execution_unit_0_alu_0_n_46_0),.B2(execution_unit_0_alu_0_n_108),.ZN(execution_unit_0_alu_0_n_46_2));
	INV_X1_LVT execution_unit_0alu_0i_46_3 (.A(execution_unit_0_alu_0_n_46_2),.ZN(execution_unit_0_alu_0_n_109));
	INV_X1_LVT execution_unit_0alu_0i_48_0 (.A(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_alu_0_n_48_0));
	NOR3_X1_LVT execution_unit_0alu_0i_48_1 (.A1(execution_unit_0_alu_0_n_48_0),.A2(execution_unit_0_alu_0_n_15),.A3(execution_unit_0_n_86),.ZN(execution_unit_0_alu_0_n_48_1));
	AOI21_X1_LVT execution_unit_0alu_0i_48_2 (.A(execution_unit_0_alu_0_n_48_1),.B1(execution_unit_0_alu_0_n_48_0),.B2(execution_unit_0_alu_0_n_110),.ZN(execution_unit_0_alu_0_n_48_2));
	INV_X1_LVT execution_unit_0alu_0i_48_3 (.A(execution_unit_0_alu_0_n_48_2),.ZN(execution_unit_0_alu_0_n_111));
	AOI22_X1_LVT execution_unit_0alu_0i_51_25 (.A1(execution_unit_0_alu_0_n_51_8),.A2(execution_unit_0_alu_0_n_109),.B1(inst_bw),.B2(execution_unit_0_alu_0_n_111),.ZN(execution_unit_0_alu_0_n_51_22));
	OAI22_X1_LVT execution_unit_0alu_0i_51_26 (.A1(execution_unit_0_alu_0_n_51_2),.A2(execution_unit_0_alu_0_n_51_21),.B1(execution_unit_0_alu_0_n_51_7),.B2(execution_unit_0_alu_0_n_51_22),.ZN(execution_unit_0_alu_stat[3]));
	INV_X1_LVT execution_unit_0alu_0i_51_21 (.A(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_alu_0_n_51_19));
	INV_X1_LVT execution_unit_0alu_0i_51_22 (.A(execution_unit_0_alu_out[15]),.ZN(execution_unit_0_alu_0_n_51_20));
	OAI22_X1_LVT execution_unit_0alu_0i_51_23 (.A1(execution_unit_0_alu_0_n_51_8),.A2(execution_unit_0_alu_0_n_51_19),.B1(execution_unit_0_alu_0_n_51_20),.B2(inst_bw),.ZN(execution_unit_0_alu_stat[2]));
	OR4_X1_LVT execution_unit_0alu_0i_51_11 (.A1(execution_unit_0_alu_0_n_51_8),.A2(execution_unit_0_alu_out[5]),.A3(execution_unit_0_alu_out[6]),.A4(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_alu_0_n_51_10));
	OR4_X1_LVT execution_unit_0alu_0i_51_12 (.A1(execution_unit_0_alu_0_n_51_10),.A2(execution_unit_0_alu_out[2]),.A3(execution_unit_0_alu_out[3]),.A4(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_alu_0_n_51_11));
	OR3_X1_LVT execution_unit_0alu_0i_51_13 (.A1(execution_unit_0_alu_0_n_51_11),.A2(execution_unit_0_alu_out[0]),.A3(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_alu_0_n_51_12));
	NOR4_X1_LVT execution_unit_0alu_0i_51_14 (.A1(execution_unit_0_alu_out[13]),.A2(execution_unit_0_alu_out[14]),.A3(execution_unit_0_alu_out[15]),.A4(inst_bw),.ZN(execution_unit_0_alu_0_n_51_13));
	NOR4_X1_LVT execution_unit_0alu_0i_51_15 (.A1(execution_unit_0_alu_out[4]),.A2(execution_unit_0_alu_out[5]),.A3(execution_unit_0_alu_out[6]),.A4(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_alu_0_n_51_14));
	NOR4_X1_LVT execution_unit_0alu_0i_51_16 (.A1(execution_unit_0_alu_out[9]),.A2(execution_unit_0_alu_out[10]),.A3(execution_unit_0_alu_out[11]),.A4(execution_unit_0_alu_out[12]),.ZN(execution_unit_0_alu_0_n_51_15));
	INV_X1_LVT execution_unit_0alu_0i_51_17 (.A(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_alu_0_n_51_16));
	NAND4_X1_LVT execution_unit_0alu_0i_51_18 (.A1(execution_unit_0_alu_0_n_51_13),.A2(execution_unit_0_alu_0_n_51_14),.A3(execution_unit_0_alu_0_n_51_15),.A4(execution_unit_0_alu_0_n_51_16),.ZN(execution_unit_0_alu_0_n_51_17));
	OR4_X1_LVT execution_unit_0alu_0i_51_19 (.A1(execution_unit_0_alu_0_n_51_17),.A2(execution_unit_0_alu_out[0]),.A3(execution_unit_0_alu_out[1]),.A4(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_alu_0_n_51_18));
	OAI21_X1_LVT execution_unit_0alu_0i_51_20 (.A(execution_unit_0_alu_0_n_51_12),.B1(execution_unit_0_alu_0_n_51_18),.B2(execution_unit_0_alu_out[8]),.ZN(execution_unit_0_alu_stat[1]));
	NAND2_X1_LVT execution_unit_0alu_0i_51_0 (.A1(execution_unit_0_alu_0_n_8),.A2(inst_alu[10]),.ZN(execution_unit_0_alu_0_n_51_0));
	INV_X1_LVT execution_unit_0alu_0i_51_3 (.A(inst_alu[8]),.ZN(execution_unit_0_alu_0_n_51_3));
	OAI21_X1_LVT execution_unit_0alu_0i_51_4 (.A(execution_unit_0_alu_0_n_51_2),.B1(inst_alu[10]),.B2(execution_unit_0_alu_0_n_51_3),.ZN(execution_unit_0_alu_0_n_51_4));
	INV_X1_LVT execution_unit_0alu_0i_49_0 (.A(inst_bw),.ZN(execution_unit_0_alu_0_n_49_0));
	OR4_X1_LVT execution_unit_0alu_0i_49_1 (.A1(execution_unit_0_alu_0_n_49_0),.A2(execution_unit_0_alu_out[5]),.A3(execution_unit_0_alu_out[6]),.A4(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_alu_0_n_49_1));
	OR4_X1_LVT execution_unit_0alu_0i_49_2 (.A1(execution_unit_0_alu_0_n_49_1),.A2(execution_unit_0_alu_out[2]),.A3(execution_unit_0_alu_out[3]),.A4(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_alu_0_n_49_2));
	OR3_X1_LVT execution_unit_0alu_0i_49_3 (.A1(execution_unit_0_alu_0_n_49_2),.A2(execution_unit_0_alu_out[0]),.A3(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_alu_0_n_49_3));
	NOR4_X1_LVT execution_unit_0alu_0i_49_4 (.A1(execution_unit_0_alu_out[13]),.A2(execution_unit_0_alu_out[14]),.A3(execution_unit_0_alu_out[15]),.A4(inst_bw),.ZN(execution_unit_0_alu_0_n_49_4));
	NOR4_X1_LVT execution_unit_0alu_0i_49_5 (.A1(execution_unit_0_alu_out[5]),.A2(execution_unit_0_alu_out[6]),.A3(execution_unit_0_alu_out[7]),.A4(execution_unit_0_alu_out[8]),.ZN(execution_unit_0_alu_0_n_49_5));
	NOR4_X1_LVT execution_unit_0alu_0i_49_6 (.A1(execution_unit_0_alu_out[9]),.A2(execution_unit_0_alu_out[10]),.A3(execution_unit_0_alu_out[11]),.A4(execution_unit_0_alu_out[12]),.ZN(execution_unit_0_alu_0_n_49_6));
	INV_X1_LVT execution_unit_0alu_0i_49_7 (.A(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_alu_0_n_49_7));
	NAND4_X1_LVT execution_unit_0alu_0i_49_8 (.A1(execution_unit_0_alu_0_n_49_4),.A2(execution_unit_0_alu_0_n_49_5),.A3(execution_unit_0_alu_0_n_49_6),.A4(execution_unit_0_alu_0_n_49_7),.ZN(execution_unit_0_alu_0_n_49_8));
	OR4_X1_LVT execution_unit_0alu_0i_49_9 (.A1(execution_unit_0_alu_0_n_49_8),.A2(execution_unit_0_alu_out[1]),.A3(execution_unit_0_alu_out[2]),.A4(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_alu_0_n_49_9));
	OAI21_X1_LVT execution_unit_0alu_0i_49_10 (.A(execution_unit_0_alu_0_n_49_3),.B1(execution_unit_0_alu_0_n_49_9),.B2(execution_unit_0_alu_out[0]),.ZN(execution_unit_0_alu_0_Z));
	INV_X1_LVT execution_unit_0alu_0i_50_0 (.A(execution_unit_0_alu_0_Z),.ZN(execution_unit_0_alu_0_n_112));
	NAND2_X1_LVT execution_unit_0alu_0i_51_5 (.A1(execution_unit_0_alu_0_n_51_4),.A2(execution_unit_0_alu_0_n_112),.ZN(execution_unit_0_alu_0_n_51_5));
	XNOR2_X1_LVT execution_unit_0alu_0i_41_16 (.A(execution_unit_0_alu_0_alu_add[0]),.B(execution_unit_0_alu_0_n_41_15),.ZN(execution_unit_0_alu_0_n_41_16));
	INV_X1_LVT execution_unit_0alu_0i_41_17 (.A(execution_unit_0_alu_0_n_41_16),.ZN(execution_unit_0_alu_0_alu_add_inc[0]));
	OR2_X1_LVT execution_unit_0alu_0i_27_7 (.A1(execution_unit_0_alu_0_n_82),.A2(execution_unit_0_alu_0_n_84),.ZN(execution_unit_0_alu_0_n_27_5));
	HA_X1_LVT execution_unit_0alu_0i_26_2 (.A(execution_unit_0_alu_0_n_80),.B(execution_unit_0_alu_0_n_26_1),.CO(execution_unit_0_alu_0_n_26_2),.S(execution_unit_0_alu_0_n_85));
	INV_X1_LVT execution_unit_0alu_0i_27_8 (.A(execution_unit_0_alu_0_n_85),.ZN(execution_unit_0_alu_0_n_27_6));
	XNOR2_X1_LVT execution_unit_0alu_0i_27_10 (.A(execution_unit_0_alu_0_n_27_5),.B(execution_unit_0_alu_0_n_27_6),.ZN(execution_unit_0_alu_0_n_27_8));
	XNOR2_X1_LVT execution_unit_0alu_0i_27_11 (.A(execution_unit_0_alu_0_n_27_8),.B(execution_unit_0_alu_0_n_27_7),.ZN(execution_unit_0_alu_0_bcd_add2[4]));
	AOI22_X1_LVT execution_unit_0alu_0i_44_32 (.A1(execution_unit_0_alu_0_n_104),.A2(execution_unit_0_alu_0_alu_add_inc[0]),.B1(execution_unit_0_alu_0_n_106),.B2(execution_unit_0_alu_0_bcd_add2[4]),.ZN(execution_unit_0_alu_0_n_44_16));
	INV_X1_LVT execution_unit_0alu_0i_44_33 (.A(execution_unit_0_alu_0_n_44_16),.ZN(execution_unit_0_alu_0_n_107));
	AOI22_X1_LVT execution_unit_0alu_0i_51_9 (.A1(execution_unit_0_alu_0_n_51_8),.A2(execution_unit_0_alu_0_n_107),.B1(execution_unit_0_alu_out[8]),.B2(inst_bw),.ZN(execution_unit_0_alu_0_n_51_9));
	OAI211_X1_LVT execution_unit_0alu_0i_51_10 (.A(execution_unit_0_alu_0_n_51_0),.B(execution_unit_0_alu_0_n_51_5),.C1(execution_unit_0_alu_0_n_51_7),.C2(execution_unit_0_alu_0_n_51_9),.ZN(execution_unit_0_alu_stat[0]));
	AND2_X1_LVT execution_unit_0alu_0i_52_0 (.A1(inst_alu[9]),.A2(execution_unit_0_n_0),.ZN(execution_unit_0_alu_stat_wr[0]));
	NAND3_X1_LVT execution_unit_0i_21_0 (.A1(inst_type[2]),.A2(inst_ad[0]),.A3(execution_unit_0_n_13),.ZN(execution_unit_0_n_21_0));
	NAND3_X1_LVT execution_unit_0i_21_1 (.A1(inst_as[0]),.A2(execution_unit_0_n_39),.A3(inst_type[0]),.ZN(execution_unit_0_n_21_1));
	INV_X1_LVT execution_unit_0i_21_2 (.A(inst_type[1]),.ZN(execution_unit_0_n_21_2));
	NAND3_X1_LVT execution_unit_0i_21_3 (.A1(execution_unit_0_n_21_0),.A2(execution_unit_0_n_21_1),.A3(execution_unit_0_n_21_2),.ZN(execution_unit_0_n_21_3));
	AOI21_X1_LVT execution_unit_0i_21_4 (.A(dbg_reg_wr),.B1(execution_unit_0_n_21_3),.B2(execution_unit_0_n_0),.ZN(execution_unit_0_n_21_4));
	INV_X1_LVT execution_unit_0i_21_5 (.A(execution_unit_0_n_21_4),.ZN(execution_unit_0_reg_dest_wr));
	AOI21_X1_LVT execution_unit_0i_23_0 (.A(execution_unit_0_n_40),.B1(inst_so[5]),.B2(execution_unit_0_n_0),.ZN(execution_unit_0_n_23_0));
	INV_X1_LVT execution_unit_0i_23_1 (.A(execution_unit_0_n_23_0),.ZN(execution_unit_0_reg_pc_call));
	AND2_X1_LVT execution_unit_0i_30_0 (.A1(execution_unit_0_n_11),.A2(execution_unit_0_n_46),.ZN(execution_unit_0_n_30_0));
	INV_X1_LVT execution_unit_0i_30_1 (.A(execution_unit_0_n_45),.ZN(execution_unit_0_n_30_1));
	NOR3_X1_LVT execution_unit_0i_30_2 (.A1(execution_unit_0_n_30_1),.A2(execution_unit_0_n_42),.A3(inst_as[1]),.ZN(execution_unit_0_n_30_2));
	OR4_X1_LVT execution_unit_0i_30_3 (.A1(execution_unit_0_n_30_0),.A2(execution_unit_0_n_30_2),.A3(execution_unit_0_n_44),.A4(execution_unit_0_n_43),.ZN(execution_unit_0_reg_sp_wr));
	AOI221_X1_LVT execution_unit_0i_32_0 (.A(execution_unit_0_n_9),.B1(exec_done),.B2(inst_as[3]),.C1(execution_unit_0_n_1),.C2(inst_so[6]),.ZN(execution_unit_0_n_32_0));
	INV_X1_LVT execution_unit_0i_32_1 (.A(execution_unit_0_n_32_0),.ZN(execution_unit_0_reg_incr));
	INV_X1_LVT execution_unit_0register_file_0i_6_0 (.A(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_6_0));
	AOI21_X1_LVT execution_unit_0register_file_0i_1_0 (.A(execution_unit_0_reg_sr_wr),.B1(inst_dest[2]),.B2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_n_1_0));
	INV_X1_LVT execution_unit_0register_file_0i_1_1 (.A(execution_unit_0_register_file_0_n_1_0),.ZN(execution_unit_0_register_file_0_r2_wr));
	INV_X1_LVT execution_unit_0register_file_0i_2_0 (.A(execution_unit_0_register_file_0_r2_wr),.ZN(execution_unit_0_register_file_0_n_2_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_2_3 (.A1(execution_unit_0_register_file_0_n_2_0),.A2(execution_unit_0_register_file_0_n_7),.B1(execution_unit_0_register_file_0_r2_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_2_2));
	INV_X1_LVT execution_unit_0register_file_0i_2_4 (.A(execution_unit_0_register_file_0_n_2_2),.ZN(execution_unit_0_register_file_0_r2_nxt[1]));
	AND2_X1_LVT execution_unit_0register_file_0i_6_5 (.A1(execution_unit_0_register_file_0_n_6_0),.A2(execution_unit_0_register_file_0_r2_nxt[1]),.ZN(execution_unit_0_register_file_0_n_17));
	INV_X1_LVT execution_unit_0register_file_0i_3_0 (.A(puc_rst),.ZN(execution_unit_0_register_file_0_n_8));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_17),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_register_file_0_n_7),.QN());
	AOI21_X1_LVT execution_unit_0register_file_0i_8_0 (.A(execution_unit_0_register_file_0_n_7),.B1(execution_unit_0_register_file_0_r2_nxt[1]),.B2(execution_unit_0_register_file_0_r2_wr),.ZN(execution_unit_0_register_file_0_n_8_0));
	INV_X1_LVT execution_unit_0register_file_0i_8_1 (.A(execution_unit_0_register_file_0_n_8_0),.ZN(cpuoff));
	AOI22_X1_LVT execution_unit_0register_file_0i_2_1 (.A1(execution_unit_0_register_file_0_n_2_0),.A2(gie),.B1(execution_unit_0_alu_out[3]),.B2(execution_unit_0_register_file_0_r2_wr),.ZN(execution_unit_0_register_file_0_n_2_1));
	INV_X1_LVT execution_unit_0register_file_0i_2_2 (.A(execution_unit_0_register_file_0_n_2_1),.ZN(execution_unit_0_register_file_0_r2_nxt[0]));
	AND2_X1_LVT execution_unit_0register_file_0i_6_4 (.A1(execution_unit_0_register_file_0_n_6_0),.A2(execution_unit_0_register_file_0_r2_nxt[0]),.ZN(execution_unit_0_register_file_0_n_16));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_16),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(gie),.QN());
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b5___05F05d (.D(1'b0),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(oscoff),.QN());
	INV_X1_LVT execution_unit_0register_file_0i_0_0 (.A(inst_bw),.ZN(execution_unit_0_register_file_0_n_0_0));
	AND2_X1_LVT execution_unit_0register_file_0i_0_8 (.A1(execution_unit_0_register_file_0_n_0_0),.A2(execution_unit_0_alu_out[15]),.ZN(pc_sw[15]));
	AND2_X1_LVT execution_unit_0register_file_0i_0_7 (.A1(execution_unit_0_register_file_0_n_0_0),.A2(execution_unit_0_alu_out[14]),.ZN(pc_sw[14]));
	AND2_X1_LVT execution_unit_0register_file_0i_0_6 (.A1(execution_unit_0_register_file_0_n_0_0),.A2(execution_unit_0_alu_out[13]),.ZN(pc_sw[13]));
	AND2_X1_LVT execution_unit_0register_file_0i_0_5 (.A1(execution_unit_0_register_file_0_n_0_0),.A2(execution_unit_0_alu_out[12]),.ZN(pc_sw[12]));
	AND2_X1_LVT execution_unit_0register_file_0i_0_4 (.A1(execution_unit_0_register_file_0_n_0_0),.A2(execution_unit_0_alu_out[11]),.ZN(pc_sw[11]));
	AND2_X1_LVT execution_unit_0register_file_0i_0_3 (.A1(execution_unit_0_register_file_0_n_0_0),.A2(execution_unit_0_alu_out[10]),.ZN(pc_sw[10]));
	AND2_X1_LVT execution_unit_0register_file_0i_0_2 (.A1(execution_unit_0_register_file_0_n_0_0),.A2(execution_unit_0_alu_out[9]),.ZN(pc_sw[9]));
	AND2_X1_LVT execution_unit_0register_file_0i_0_1 (.A1(execution_unit_0_register_file_0_n_0_0),.A2(execution_unit_0_alu_out[8]),.ZN(pc_sw[8]));
	AOI21_X1_LVT execution_unit_0register_file_0i_9_0 (.A(execution_unit_0_reg_pc_call),.B1(inst_dest[0]),.B2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_n_9_0));
	INV_X1_LVT execution_unit_0register_file_0i_9_1 (.A(execution_unit_0_register_file_0_n_9_0),.ZN(pc_sw_wr));
	AND2_X1_LVT execution_unit_0register_file_0i_19_0 (.A1(inst_dest[4]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r4_wr));
	INV_X1_LVT execution_unit_0register_file_0i_24_0 (.A(execution_unit_0_register_file_0_r4_wr),.ZN(execution_unit_0_register_file_0_n_24_0));
	INV_X1_LVT execution_unit_0register_file_0i_17_0 (.A(inst_src[4]),.ZN(execution_unit_0_register_file_0_n_17_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_17_1 (.A1(execution_unit_0_register_file_0_n_17_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_24));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_315 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[15]),.ZN(execution_unit_0_register_file_0_n_105_300));
	INV_X1_LVT execution_unit_0register_file_0i_14_0 (.A(inst_src[3]),.ZN(execution_unit_0_register_file_0_n_14_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_14_1 (.A1(execution_unit_0_register_file_0_n_14_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_22));
	AND2_X1_LVT execution_unit_0register_file_0i_15_0 (.A1(inst_dest[3]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r3_wr));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r3_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_r3_wr),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_23));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b15___05F05d (.D(pc_sw[15]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_316 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[15]),.ZN(execution_unit_0_register_file_0_n_105_301));
	INV_X1_LVT execution_unit_0register_file_0i_13_1 (.A(inst_src[2]),.ZN(execution_unit_0_register_file_0_n_13_1));
	INV_X1_LVT execution_unit_0register_file_0i_13_0 (.A(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_13_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_13_2 (.A1(execution_unit_0_register_file_0_n_13_1),.A2(execution_unit_0_register_file_0_n_13_0),.ZN(execution_unit_0_register_file_0_n_21));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b15___05F05d (.D(1'b0),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_register_file_0_n_0),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_317 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_register_file_0_n_0),.ZN(execution_unit_0_register_file_0_n_105_302));
	INV_X1_LVT execution_unit_0register_file_0i_10_0 (.A(inst_src[1]),.ZN(execution_unit_0_register_file_0_n_10_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_10_1 (.A1(execution_unit_0_register_file_0_n_10_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_inst_src_in));
	AND2_X1_LVT execution_unit_0register_file_0i_12_0 (.A1(inst_dest[1]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r1_wr));
	INV_X1_LVT execution_unit_0register_file_0i_108_1 (.A(execution_unit_0_reg_sp_wr),.ZN(execution_unit_0_register_file_0_n_108_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_108_2 (.A1(execution_unit_0_register_file_0_n_108_0),.A2(execution_unit_0_register_file_0_r1_wr),.ZN(execution_unit_0_register_file_0_n_272));
	NOR2_X1_LVT execution_unit_0register_file_0i_108_0 (.A1(execution_unit_0_reg_sp_wr),.A2(execution_unit_0_register_file_0_r1_wr),.ZN(execution_unit_0_register_file_0_n_271));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_27 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_24_14));
	INV_X1_LVT execution_unit_0register_file_0i_24_28 (.A(execution_unit_0_register_file_0_n_24_14),.ZN(execution_unit_0_register_file_0_n_41));
	AND2_X1_LVT execution_unit_0register_file_0i_18_0 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r4_inc));
	INV_X1_LVT execution_unit_0register_file_0i_25_1 (.A(execution_unit_0_register_file_0_r4_inc),.ZN(execution_unit_0_register_file_0_n_25_1));
	INV_X1_LVT execution_unit_0register_file_0i_25_0 (.A(execution_unit_0_register_file_0_r4_wr),.ZN(execution_unit_0_register_file_0_n_25_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_25_2 (.A1(execution_unit_0_register_file_0_n_25_1),.A2(execution_unit_0_register_file_0_n_25_0),.ZN(execution_unit_0_register_file_0_n_44));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r4_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_44),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_27));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_41),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_273 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[13]),.ZN(execution_unit_0_register_file_0_n_105_260));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b13___05F05d (.D(pc_sw[13]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_274 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[13]),.ZN(execution_unit_0_register_file_0_n_105_261));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b13___05F05d (.D(1'b0),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_register_file_0_n_2),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_275 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_register_file_0_n_2),.ZN(execution_unit_0_register_file_0_n_105_262));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_23 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_24_12));
	INV_X1_LVT execution_unit_0register_file_0i_24_24 (.A(execution_unit_0_register_file_0_n_24_12),.ZN(execution_unit_0_register_file_0_n_39));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_39),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_231 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[11]),.ZN(execution_unit_0_register_file_0_n_105_220));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b11___05F05d (.D(pc_sw[11]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_232 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[11]),.ZN(execution_unit_0_register_file_0_n_105_221));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b11___05F05d (.D(1'b0),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_register_file_0_n_4),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_233 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_register_file_0_n_4),.ZN(execution_unit_0_register_file_0_n_105_222));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_19 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_24_10));
	INV_X1_LVT execution_unit_0register_file_0i_24_20 (.A(execution_unit_0_register_file_0_n_24_10),.ZN(execution_unit_0_register_file_0_n_37));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_37),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_189 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[9]),.ZN(execution_unit_0_register_file_0_n_105_180));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b9___05F05d (.D(pc_sw[9]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_190 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[9]),.ZN(execution_unit_0_register_file_0_n_105_181));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b9___05F05d (.D(1'b0),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_register_file_0_n_6),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_191 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_register_file_0_n_6),.ZN(execution_unit_0_register_file_0_n_105_182));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_15 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_24_8));
	INV_X1_LVT execution_unit_0register_file_0i_24_16 (.A(execution_unit_0_register_file_0_n_24_8),.ZN(execution_unit_0_register_file_0_n_35));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_35),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_147 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[7]),.ZN(execution_unit_0_register_file_0_n_105_140));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b7___05F05d (.D(execution_unit_0_alu_out[7]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_148 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[7]),.ZN(execution_unit_0_register_file_0_n_105_141));
	AOI22_X1_LVT execution_unit_0register_file_0i_2_7 (.A1(execution_unit_0_register_file_0_n_2_0),.A2(scg1),.B1(execution_unit_0_register_file_0_r2_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_2_4));
	INV_X1_LVT execution_unit_0register_file_0i_2_8 (.A(execution_unit_0_register_file_0_n_2_4),.ZN(execution_unit_0_register_file_0_r2_nxt[4]));
	AND2_X1_LVT execution_unit_0register_file_0i_6_7 (.A1(execution_unit_0_register_file_0_n_6_0),.A2(execution_unit_0_register_file_0_r2_nxt[4]),.ZN(execution_unit_0_register_file_0_n_19));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_19),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(scg1),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_149 (.A1(execution_unit_0_register_file_0_n_21),.A2(scg1),.ZN(execution_unit_0_register_file_0_n_105_142));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_11 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_24_6));
	INV_X1_LVT execution_unit_0register_file_0i_24_12 (.A(execution_unit_0_register_file_0_n_24_6),.ZN(execution_unit_0_register_file_0_n_33));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_33),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_105 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[5]),.ZN(execution_unit_0_register_file_0_n_105_100));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b5___05F05d (.D(execution_unit_0_alu_out[5]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_106 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[5]),.ZN(execution_unit_0_register_file_0_n_105_101));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_107 (.A1(execution_unit_0_register_file_0_n_21),.A2(oscoff),.ZN(execution_unit_0_register_file_0_n_105_102));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_7 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_24_4));
	INV_X1_LVT execution_unit_0register_file_0i_24_8 (.A(execution_unit_0_register_file_0_n_24_4),.ZN(execution_unit_0_register_file_0_n_31));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_31),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_63 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[3]),.ZN(execution_unit_0_register_file_0_n_105_60));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b3___05F05d (.D(execution_unit_0_alu_out[3]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_64 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[3]),.ZN(execution_unit_0_register_file_0_n_105_61));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_65 (.A1(execution_unit_0_register_file_0_n_21),.A2(gie),.ZN(execution_unit_0_register_file_0_n_105_62));
	INV_X1_LVT execution_unit_0register_file_0i_20_0 (.A(inst_bw),.ZN(execution_unit_0_register_file_0_n_20_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_20_1 (.A1(execution_unit_0_register_file_0_n_20_0),.A2(execution_unit_0_register_file_0_inst_src_in),.ZN(execution_unit_0_register_file_0_n_25));
	INV_X1_LVT execution_unit_0register_file_0i_21_0 (.A(execution_unit_0_register_file_0_n_25),.ZN(execution_unit_0_register_file_0_n_26));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_3 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_24_2));
	INV_X1_LVT execution_unit_0register_file_0i_24_4 (.A(execution_unit_0_register_file_0_n_24_2),.ZN(execution_unit_0_register_file_0_n_29));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_29),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_21 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[1]),.ZN(execution_unit_0_register_file_0_n_105_20));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b1___05F05d (.D(execution_unit_0_alu_out[1]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_22 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[1]),.ZN(execution_unit_0_register_file_0_n_105_21));
	INV_X1_LVT execution_unit_0register_file_0i_5_0 (.A(execution_unit_0_register_file_0_r2_wr),.ZN(execution_unit_0_register_file_0_n_5_0));
	INV_X1_LVT execution_unit_0register_file_0i_5_6 (.A(execution_unit_0_alu_stat_wr[1]),.ZN(execution_unit_0_register_file_0_n_5_5));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_7 (.A1(execution_unit_0_register_file_0_n_5_0),.A2(execution_unit_0_register_file_0_n_5_5),.A3(execution_unit_0_status[1]),.ZN(execution_unit_0_register_file_0_n_5_6));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_8 (.A1(execution_unit_0_register_file_0_n_5_5),.A2(execution_unit_0_register_file_0_r2_wr),.A3(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_5_7));
	NAND2_X1_LVT execution_unit_0register_file_0i_5_9 (.A1(execution_unit_0_alu_stat[1]),.A2(execution_unit_0_alu_stat_wr[1]),.ZN(execution_unit_0_register_file_0_n_5_8));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_10 (.A1(execution_unit_0_register_file_0_n_5_6),.A2(execution_unit_0_register_file_0_n_5_7),.A3(execution_unit_0_register_file_0_n_5_8),.ZN(execution_unit_0_register_file_0_n_10));
	AND2_X1_LVT execution_unit_0register_file_0i_6_2 (.A1(execution_unit_0_register_file_0_n_6_0),.A2(execution_unit_0_register_file_0_n_10),.ZN(execution_unit_0_register_file_0_n_14));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_14),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_status[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_23 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_status[1]),.ZN(execution_unit_0_register_file_0_n_105_22));
	INV_X1_LVT execution_unit_0register_file_0i_106_0 (.A(execution_unit_0_reg_src[1]),.ZN(execution_unit_0_register_file_0_n_255));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_0 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(execution_unit_0_alu_out[1]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[1]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_255),.ZN(execution_unit_0_register_file_0_n_109_0));
	INV_X1_LVT execution_unit_0register_file_0i_109_1 (.A(execution_unit_0_register_file_0_n_109_0),.ZN(execution_unit_0_register_file_0_n_273));
	INV_X1_LVT execution_unit_0register_file_0i_110_0 (.A(execution_unit_0_reg_sp_wr),.ZN(execution_unit_0_register_file_0_n_110_0));
	INV_X1_LVT execution_unit_0register_file_0i_110_1 (.A(execution_unit_0_register_file_0_r1_wr),.ZN(execution_unit_0_register_file_0_n_110_1));
	AND2_X1_LVT execution_unit_0register_file_0i_11_0 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r1_inc));
	NAND3_X1_LVT execution_unit_0register_file_0i_110_2 (.A1(execution_unit_0_register_file_0_n_110_0),.A2(execution_unit_0_register_file_0_n_110_1),.A3(execution_unit_0_register_file_0_r1_inc),.ZN(execution_unit_0_register_file_0_n_110_2));
	NAND3_X1_LVT execution_unit_0register_file_0i_110_3 (.A1(execution_unit_0_register_file_0_n_110_2),.A2(execution_unit_0_register_file_0_n_110_0),.A3(execution_unit_0_register_file_0_n_110_1),.ZN(execution_unit_0_register_file_0_n_288));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r1_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_288),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_270));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_273),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_24 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[1]),.ZN(execution_unit_0_register_file_0_n_105_23));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_25 (.A1(execution_unit_0_register_file_0_n_105_20),.A2(execution_unit_0_register_file_0_n_105_21),.A3(execution_unit_0_register_file_0_n_105_22),.A4(execution_unit_0_register_file_0_n_105_23),.ZN(execution_unit_0_register_file_0_n_105_24));
	INV_X1_LVT execution_unit_0register_file_0i_76_0 (.A(inst_src[12]),.ZN(execution_unit_0_register_file_0_n_76_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_76_1 (.A1(execution_unit_0_register_file_0_n_76_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_178));
	AND2_X1_LVT execution_unit_0register_file_0i_78_0 (.A1(inst_dest[12]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r12_wr));
	INV_X1_LVT execution_unit_0register_file_0i_80_0 (.A(execution_unit_0_register_file_0_r12_wr),.ZN(execution_unit_0_register_file_0_n_80_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_3 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_80_2));
	INV_X1_LVT execution_unit_0register_file_0i_80_4 (.A(execution_unit_0_register_file_0_n_80_2),.ZN(execution_unit_0_register_file_0_n_181));
	AND2_X1_LVT execution_unit_0register_file_0i_77_0 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r12_inc));
	INV_X1_LVT execution_unit_0register_file_0i_81_1 (.A(execution_unit_0_register_file_0_r12_inc),.ZN(execution_unit_0_register_file_0_n_81_1));
	INV_X1_LVT execution_unit_0register_file_0i_81_0 (.A(execution_unit_0_register_file_0_r12_wr),.ZN(execution_unit_0_register_file_0_n_81_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_81_2 (.A1(execution_unit_0_register_file_0_n_81_1),.A2(execution_unit_0_register_file_0_n_81_0),.ZN(execution_unit_0_register_file_0_n_196));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r12_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_196),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_179));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_181),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_26 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[1]),.ZN(execution_unit_0_register_file_0_n_105_25));
	INV_X1_LVT execution_unit_0register_file_0i_69_0 (.A(inst_src[11]),.ZN(execution_unit_0_register_file_0_n_69_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_69_1 (.A1(execution_unit_0_register_file_0_n_69_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_159));
	AND2_X1_LVT execution_unit_0register_file_0i_71_0 (.A1(inst_dest[11]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r11_wr));
	INV_X1_LVT execution_unit_0register_file_0i_73_0 (.A(execution_unit_0_register_file_0_r11_wr),.ZN(execution_unit_0_register_file_0_n_73_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_3 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_73_2));
	INV_X1_LVT execution_unit_0register_file_0i_73_4 (.A(execution_unit_0_register_file_0_n_73_2),.ZN(execution_unit_0_register_file_0_n_162));
	AND2_X1_LVT execution_unit_0register_file_0i_70_0 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r11_inc));
	INV_X1_LVT execution_unit_0register_file_0i_74_1 (.A(execution_unit_0_register_file_0_r11_inc),.ZN(execution_unit_0_register_file_0_n_74_1));
	INV_X1_LVT execution_unit_0register_file_0i_74_0 (.A(execution_unit_0_register_file_0_r11_wr),.ZN(execution_unit_0_register_file_0_n_74_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_74_2 (.A1(execution_unit_0_register_file_0_n_74_1),.A2(execution_unit_0_register_file_0_n_74_0),.ZN(execution_unit_0_register_file_0_n_177));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r11_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_177),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_160));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_162),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_27 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[1]),.ZN(execution_unit_0_register_file_0_n_105_26));
	INV_X1_LVT execution_unit_0register_file_0i_62_0 (.A(inst_src[10]),.ZN(execution_unit_0_register_file_0_n_62_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_62_1 (.A1(execution_unit_0_register_file_0_n_62_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_140));
	AND2_X1_LVT execution_unit_0register_file_0i_64_0 (.A1(inst_dest[10]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r10_wr));
	INV_X1_LVT execution_unit_0register_file_0i_66_0 (.A(execution_unit_0_register_file_0_r10_wr),.ZN(execution_unit_0_register_file_0_n_66_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_3 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_66_2));
	INV_X1_LVT execution_unit_0register_file_0i_66_4 (.A(execution_unit_0_register_file_0_n_66_2),.ZN(execution_unit_0_register_file_0_n_143));
	AND2_X1_LVT execution_unit_0register_file_0i_63_0 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r10_inc));
	INV_X1_LVT execution_unit_0register_file_0i_67_1 (.A(execution_unit_0_register_file_0_r10_inc),.ZN(execution_unit_0_register_file_0_n_67_1));
	INV_X1_LVT execution_unit_0register_file_0i_67_0 (.A(execution_unit_0_register_file_0_r10_wr),.ZN(execution_unit_0_register_file_0_n_67_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_67_2 (.A1(execution_unit_0_register_file_0_n_67_1),.A2(execution_unit_0_register_file_0_n_67_0),.ZN(execution_unit_0_register_file_0_n_158));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r10_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_158),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_141));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_143),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_28 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[1]),.ZN(execution_unit_0_register_file_0_n_105_27));
	INV_X1_LVT execution_unit_0register_file_0i_55_0 (.A(inst_src[9]),.ZN(execution_unit_0_register_file_0_n_55_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_55_1 (.A1(execution_unit_0_register_file_0_n_55_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_121));
	AND2_X1_LVT execution_unit_0register_file_0i_57_0 (.A1(inst_dest[9]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r9_wr));
	INV_X1_LVT execution_unit_0register_file_0i_59_0 (.A(execution_unit_0_register_file_0_r9_wr),.ZN(execution_unit_0_register_file_0_n_59_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_3 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_59_2));
	INV_X1_LVT execution_unit_0register_file_0i_59_4 (.A(execution_unit_0_register_file_0_n_59_2),.ZN(execution_unit_0_register_file_0_n_124));
	AND2_X1_LVT execution_unit_0register_file_0i_56_0 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r9_inc));
	INV_X1_LVT execution_unit_0register_file_0i_60_1 (.A(execution_unit_0_register_file_0_r9_inc),.ZN(execution_unit_0_register_file_0_n_60_1));
	INV_X1_LVT execution_unit_0register_file_0i_60_0 (.A(execution_unit_0_register_file_0_r9_wr),.ZN(execution_unit_0_register_file_0_n_60_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_60_2 (.A1(execution_unit_0_register_file_0_n_60_1),.A2(execution_unit_0_register_file_0_n_60_0),.ZN(execution_unit_0_register_file_0_n_139));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r9_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_139),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_122));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_124),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_29 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[1]),.ZN(execution_unit_0_register_file_0_n_105_28));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_30 (.A1(execution_unit_0_register_file_0_n_105_25),.A2(execution_unit_0_register_file_0_n_105_26),.A3(execution_unit_0_register_file_0_n_105_27),.A4(execution_unit_0_register_file_0_n_105_28),.ZN(execution_unit_0_register_file_0_n_105_29));
	INV_X1_LVT execution_unit_0register_file_0i_48_0 (.A(inst_src[8]),.ZN(execution_unit_0_register_file_0_n_48_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_48_1 (.A1(execution_unit_0_register_file_0_n_48_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_102));
	AND2_X1_LVT execution_unit_0register_file_0i_50_0 (.A1(inst_dest[8]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r8_wr));
	INV_X1_LVT execution_unit_0register_file_0i_52_0 (.A(execution_unit_0_register_file_0_r8_wr),.ZN(execution_unit_0_register_file_0_n_52_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_3 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_52_2));
	INV_X1_LVT execution_unit_0register_file_0i_52_4 (.A(execution_unit_0_register_file_0_n_52_2),.ZN(execution_unit_0_register_file_0_n_105));
	AND2_X1_LVT execution_unit_0register_file_0i_49_0 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r8_inc));
	INV_X1_LVT execution_unit_0register_file_0i_53_1 (.A(execution_unit_0_register_file_0_r8_inc),.ZN(execution_unit_0_register_file_0_n_53_1));
	INV_X1_LVT execution_unit_0register_file_0i_53_0 (.A(execution_unit_0_register_file_0_r8_wr),.ZN(execution_unit_0_register_file_0_n_53_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_53_2 (.A1(execution_unit_0_register_file_0_n_53_1),.A2(execution_unit_0_register_file_0_n_53_0),.ZN(execution_unit_0_register_file_0_n_120));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r8_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_120),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_103));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_105),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_31 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[1]),.ZN(execution_unit_0_register_file_0_n_105_30));
	INV_X1_LVT execution_unit_0register_file_0i_41_0 (.A(inst_src[7]),.ZN(execution_unit_0_register_file_0_n_41_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_41_1 (.A1(execution_unit_0_register_file_0_n_41_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_83));
	AND2_X1_LVT execution_unit_0register_file_0i_43_0 (.A1(inst_dest[7]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r7_wr));
	INV_X1_LVT execution_unit_0register_file_0i_45_0 (.A(execution_unit_0_register_file_0_r7_wr),.ZN(execution_unit_0_register_file_0_n_45_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_3 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_45_2));
	INV_X1_LVT execution_unit_0register_file_0i_45_4 (.A(execution_unit_0_register_file_0_n_45_2),.ZN(execution_unit_0_register_file_0_n_86));
	AND2_X1_LVT execution_unit_0register_file_0i_42_0 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r7_inc));
	INV_X1_LVT execution_unit_0register_file_0i_46_1 (.A(execution_unit_0_register_file_0_r7_inc),.ZN(execution_unit_0_register_file_0_n_46_1));
	INV_X1_LVT execution_unit_0register_file_0i_46_0 (.A(execution_unit_0_register_file_0_r7_wr),.ZN(execution_unit_0_register_file_0_n_46_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_46_2 (.A1(execution_unit_0_register_file_0_n_46_1),.A2(execution_unit_0_register_file_0_n_46_0),.ZN(execution_unit_0_register_file_0_n_101));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r7_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_101),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_84));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_86),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_32 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[1]),.ZN(execution_unit_0_register_file_0_n_105_31));
	INV_X1_LVT execution_unit_0register_file_0i_34_0 (.A(inst_src[6]),.ZN(execution_unit_0_register_file_0_n_34_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_34_1 (.A1(execution_unit_0_register_file_0_n_34_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_64));
	AND2_X1_LVT execution_unit_0register_file_0i_36_0 (.A1(inst_dest[6]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r6_wr));
	INV_X1_LVT execution_unit_0register_file_0i_38_0 (.A(execution_unit_0_register_file_0_r6_wr),.ZN(execution_unit_0_register_file_0_n_38_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_3 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_38_2));
	INV_X1_LVT execution_unit_0register_file_0i_38_4 (.A(execution_unit_0_register_file_0_n_38_2),.ZN(execution_unit_0_register_file_0_n_67));
	AND2_X1_LVT execution_unit_0register_file_0i_35_0 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r6_inc));
	INV_X1_LVT execution_unit_0register_file_0i_39_1 (.A(execution_unit_0_register_file_0_r6_inc),.ZN(execution_unit_0_register_file_0_n_39_1));
	INV_X1_LVT execution_unit_0register_file_0i_39_0 (.A(execution_unit_0_register_file_0_r6_wr),.ZN(execution_unit_0_register_file_0_n_39_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_39_2 (.A1(execution_unit_0_register_file_0_n_39_1),.A2(execution_unit_0_register_file_0_n_39_0),.ZN(execution_unit_0_register_file_0_n_82));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r6_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_82),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_65));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_67),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_33 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[1]),.ZN(execution_unit_0_register_file_0_n_105_32));
	INV_X1_LVT execution_unit_0register_file_0i_27_0 (.A(inst_src[5]),.ZN(execution_unit_0_register_file_0_n_27_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_27_1 (.A1(execution_unit_0_register_file_0_n_27_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_45));
	AND2_X1_LVT execution_unit_0register_file_0i_29_0 (.A1(inst_dest[5]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r5_wr));
	INV_X1_LVT execution_unit_0register_file_0i_31_0 (.A(execution_unit_0_register_file_0_r5_wr),.ZN(execution_unit_0_register_file_0_n_31_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_3 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_31_2));
	INV_X1_LVT execution_unit_0register_file_0i_31_4 (.A(execution_unit_0_register_file_0_n_31_2),.ZN(execution_unit_0_register_file_0_n_48));
	AND2_X1_LVT execution_unit_0register_file_0i_28_0 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r5_inc));
	INV_X1_LVT execution_unit_0register_file_0i_32_1 (.A(execution_unit_0_register_file_0_r5_inc),.ZN(execution_unit_0_register_file_0_n_32_1));
	INV_X1_LVT execution_unit_0register_file_0i_32_0 (.A(execution_unit_0_register_file_0_r5_wr),.ZN(execution_unit_0_register_file_0_n_32_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_32_2 (.A1(execution_unit_0_register_file_0_n_32_1),.A2(execution_unit_0_register_file_0_n_32_0),.ZN(execution_unit_0_register_file_0_n_63));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r5_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_63),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_46));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_48),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_34 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[1]),.ZN(execution_unit_0_register_file_0_n_105_33));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_35 (.A1(execution_unit_0_register_file_0_n_105_30),.A2(execution_unit_0_register_file_0_n_105_31),.A3(execution_unit_0_register_file_0_n_105_32),.A4(execution_unit_0_register_file_0_n_105_33),.ZN(execution_unit_0_register_file_0_n_105_34));
	INV_X1_LVT execution_unit_0register_file_0i_83_0 (.A(inst_src[13]),.ZN(execution_unit_0_register_file_0_n_83_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_83_1 (.A1(execution_unit_0_register_file_0_n_83_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_197));
	AND2_X1_LVT execution_unit_0register_file_0i_85_0 (.A1(inst_dest[13]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r13_wr));
	INV_X1_LVT execution_unit_0register_file_0i_87_0 (.A(execution_unit_0_register_file_0_r13_wr),.ZN(execution_unit_0_register_file_0_n_87_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_3 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_87_2));
	INV_X1_LVT execution_unit_0register_file_0i_87_4 (.A(execution_unit_0_register_file_0_n_87_2),.ZN(execution_unit_0_register_file_0_n_200));
	AND2_X1_LVT execution_unit_0register_file_0i_84_0 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r13_inc));
	INV_X1_LVT execution_unit_0register_file_0i_88_1 (.A(execution_unit_0_register_file_0_r13_inc),.ZN(execution_unit_0_register_file_0_n_88_1));
	INV_X1_LVT execution_unit_0register_file_0i_88_0 (.A(execution_unit_0_register_file_0_r13_wr),.ZN(execution_unit_0_register_file_0_n_88_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_88_2 (.A1(execution_unit_0_register_file_0_n_88_1),.A2(execution_unit_0_register_file_0_n_88_0),.ZN(execution_unit_0_register_file_0_n_215));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r13_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_215),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_198));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_200),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[1]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_36 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[1]),.ZN(execution_unit_0_register_file_0_n_105_35));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_37 (.A1(execution_unit_0_register_file_0_n_105_24),.A2(execution_unit_0_register_file_0_n_105_29),.A3(execution_unit_0_register_file_0_n_105_34),.A4(execution_unit_0_register_file_0_n_105_35),.ZN(execution_unit_0_register_file_0_n_105_36));
	INV_X1_LVT execution_unit_0register_file_0i_104_0 (.A(inst_src[0]),.ZN(execution_unit_0_register_file_0_n_104_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_104_1 (.A1(execution_unit_0_register_file_0_n_104_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_254));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_38 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[1]),.ZN(execution_unit_0_register_file_0_n_105_37));
	INV_X1_LVT execution_unit_0register_file_0i_97_0 (.A(inst_src[15]),.ZN(execution_unit_0_register_file_0_n_97_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_97_1 (.A1(execution_unit_0_register_file_0_n_97_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_235));
	AND2_X1_LVT execution_unit_0register_file_0i_99_0 (.A1(inst_dest[15]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r15_wr));
	INV_X1_LVT execution_unit_0register_file_0i_101_0 (.A(execution_unit_0_register_file_0_r15_wr),.ZN(execution_unit_0_register_file_0_n_101_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_3 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_101_2));
	INV_X1_LVT execution_unit_0register_file_0i_101_4 (.A(execution_unit_0_register_file_0_n_101_2),.ZN(execution_unit_0_register_file_0_n_238));
	AND2_X1_LVT execution_unit_0register_file_0i_98_0 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r15_inc));
	INV_X1_LVT execution_unit_0register_file_0i_102_1 (.A(execution_unit_0_register_file_0_r15_inc),.ZN(execution_unit_0_register_file_0_n_102_1));
	INV_X1_LVT execution_unit_0register_file_0i_102_0 (.A(execution_unit_0_register_file_0_r15_wr),.ZN(execution_unit_0_register_file_0_n_102_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_102_2 (.A1(execution_unit_0_register_file_0_n_102_1),.A2(execution_unit_0_register_file_0_n_102_0),.ZN(execution_unit_0_register_file_0_n_253));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r15_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_253),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_236));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_238),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_39 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[1]),.ZN(execution_unit_0_register_file_0_n_105_38));
	INV_X1_LVT execution_unit_0register_file_0i_90_0 (.A(inst_src[14]),.ZN(execution_unit_0_register_file_0_n_90_0));
	NOR2_X1_LVT execution_unit_0register_file_0i_90_1 (.A1(execution_unit_0_register_file_0_n_90_0),.A2(execution_unit_0_reg_sr_clr),.ZN(execution_unit_0_register_file_0_n_216));
	AND2_X1_LVT execution_unit_0register_file_0i_92_0 (.A1(inst_dest[14]),.A2(execution_unit_0_reg_dest_wr),.ZN(execution_unit_0_register_file_0_r14_wr));
	INV_X1_LVT execution_unit_0register_file_0i_94_0 (.A(execution_unit_0_register_file_0_r14_wr),.ZN(execution_unit_0_register_file_0_n_94_0));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_3 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[1]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(execution_unit_0_alu_out[1]),.ZN(execution_unit_0_register_file_0_n_94_2));
	INV_X1_LVT execution_unit_0register_file_0i_94_4 (.A(execution_unit_0_register_file_0_n_94_2),.ZN(execution_unit_0_register_file_0_n_219));
	AND2_X1_LVT execution_unit_0register_file_0i_91_0 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_reg_incr),.ZN(execution_unit_0_register_file_0_r14_inc));
	INV_X1_LVT execution_unit_0register_file_0i_95_1 (.A(execution_unit_0_register_file_0_r14_inc),.ZN(execution_unit_0_register_file_0_n_95_1));
	INV_X1_LVT execution_unit_0register_file_0i_95_0 (.A(execution_unit_0_register_file_0_r14_wr),.ZN(execution_unit_0_register_file_0_n_95_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_95_2 (.A1(execution_unit_0_register_file_0_n_95_1),.A2(execution_unit_0_register_file_0_n_95_0),.ZN(execution_unit_0_register_file_0_n_234));
	CLKGATETST_X1_LVT execution_unit_0register_file_0clk_gate_r14_reg (.CK(cpu_mclk),.E(execution_unit_0_register_file_0_n_234),.SE(1'b0),.GCK(execution_unit_0_register_file_0_n_217));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b1___05F05d (.D(execution_unit_0_register_file_0_n_219),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[1]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_40 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[1]),.ZN(execution_unit_0_register_file_0_n_105_39));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_41 (.A1(execution_unit_0_register_file_0_n_105_36),.A2(execution_unit_0_register_file_0_n_105_37),.A3(execution_unit_0_register_file_0_n_105_38),.A4(execution_unit_0_register_file_0_n_105_39),.ZN(execution_unit_0_reg_src[1]));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_1 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r4_wr),.ZN(execution_unit_0_register_file_0_n_24_1));
	INV_X1_LVT execution_unit_0register_file_0i_24_2 (.A(execution_unit_0_register_file_0_n_24_1),.ZN(execution_unit_0_register_file_0_n_28));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_28),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_0 (.A1(execution_unit_0_register_file_0_r4[0]),.A2(execution_unit_0_register_file_0_n_24),.ZN(execution_unit_0_register_file_0_n_105_0));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b0___05F05d (.D(execution_unit_0_alu_out[0]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_1 (.A1(execution_unit_0_register_file_0_r3[0]),.A2(execution_unit_0_register_file_0_n_22),.ZN(execution_unit_0_register_file_0_n_105_1));
	INV_X1_LVT execution_unit_0register_file_0i_5_1 (.A(execution_unit_0_alu_stat_wr[0]),.ZN(execution_unit_0_register_file_0_n_5_1));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_2 (.A1(execution_unit_0_register_file_0_n_5_0),.A2(execution_unit_0_register_file_0_n_5_1),.A3(execution_unit_0_status[0]),.ZN(execution_unit_0_register_file_0_n_5_2));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_3 (.A1(execution_unit_0_register_file_0_n_5_1),.A2(execution_unit_0_register_file_0_r2_wr),.A3(execution_unit_0_alu_out[0]),.ZN(execution_unit_0_register_file_0_n_5_3));
	NAND2_X1_LVT execution_unit_0register_file_0i_5_4 (.A1(execution_unit_0_alu_stat[0]),.A2(execution_unit_0_alu_stat_wr[0]),.ZN(execution_unit_0_register_file_0_n_5_4));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_5 (.A1(execution_unit_0_register_file_0_n_5_2),.A2(execution_unit_0_register_file_0_n_5_3),.A3(execution_unit_0_register_file_0_n_5_4),.ZN(execution_unit_0_register_file_0_n_9));
	AND2_X1_LVT execution_unit_0register_file_0i_6_1 (.A1(execution_unit_0_register_file_0_n_6_0),.A2(execution_unit_0_register_file_0_n_9),.ZN(execution_unit_0_register_file_0_n_13));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_13),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_status[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_2 (.A1(execution_unit_0_status[0]),.A2(execution_unit_0_register_file_0_n_21),.ZN(execution_unit_0_register_file_0_n_105_2));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b0___05F05d (.D(1'b0),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_3 (.A1(execution_unit_0_register_file_0_r1[0]),.A2(execution_unit_0_register_file_0_inst_src_in),.ZN(execution_unit_0_register_file_0_n_105_3));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_4 (.A1(execution_unit_0_register_file_0_n_105_0),.A2(execution_unit_0_register_file_0_n_105_1),.A3(execution_unit_0_register_file_0_n_105_2),.A4(execution_unit_0_register_file_0_n_105_3),.ZN(execution_unit_0_register_file_0_n_105_4));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_1 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r12_wr),.ZN(execution_unit_0_register_file_0_n_80_1));
	INV_X1_LVT execution_unit_0register_file_0i_80_2 (.A(execution_unit_0_register_file_0_n_80_1),.ZN(execution_unit_0_register_file_0_n_180));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_180),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_5 (.A1(execution_unit_0_register_file_0_r12[0]),.A2(execution_unit_0_register_file_0_n_178),.ZN(execution_unit_0_register_file_0_n_105_5));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_1 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r11_wr),.ZN(execution_unit_0_register_file_0_n_73_1));
	INV_X1_LVT execution_unit_0register_file_0i_73_2 (.A(execution_unit_0_register_file_0_n_73_1),.ZN(execution_unit_0_register_file_0_n_161));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_161),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_6 (.A1(execution_unit_0_register_file_0_r11[0]),.A2(execution_unit_0_register_file_0_n_159),.ZN(execution_unit_0_register_file_0_n_105_6));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_1 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r10_wr),.ZN(execution_unit_0_register_file_0_n_66_1));
	INV_X1_LVT execution_unit_0register_file_0i_66_2 (.A(execution_unit_0_register_file_0_n_66_1),.ZN(execution_unit_0_register_file_0_n_142));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_142),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_7 (.A1(execution_unit_0_register_file_0_r10[0]),.A2(execution_unit_0_register_file_0_n_140),.ZN(execution_unit_0_register_file_0_n_105_7));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_1 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r9_wr),.ZN(execution_unit_0_register_file_0_n_59_1));
	INV_X1_LVT execution_unit_0register_file_0i_59_2 (.A(execution_unit_0_register_file_0_n_59_1),.ZN(execution_unit_0_register_file_0_n_123));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_123),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_8 (.A1(execution_unit_0_register_file_0_r9[0]),.A2(execution_unit_0_register_file_0_n_121),.ZN(execution_unit_0_register_file_0_n_105_8));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_9 (.A1(execution_unit_0_register_file_0_n_105_5),.A2(execution_unit_0_register_file_0_n_105_6),.A3(execution_unit_0_register_file_0_n_105_7),.A4(execution_unit_0_register_file_0_n_105_8),.ZN(execution_unit_0_register_file_0_n_105_9));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_1 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r8_wr),.ZN(execution_unit_0_register_file_0_n_52_1));
	INV_X1_LVT execution_unit_0register_file_0i_52_2 (.A(execution_unit_0_register_file_0_n_52_1),.ZN(execution_unit_0_register_file_0_n_104));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_104),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_10 (.A1(execution_unit_0_register_file_0_r8[0]),.A2(execution_unit_0_register_file_0_n_102),.ZN(execution_unit_0_register_file_0_n_105_10));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_1 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r7_wr),.ZN(execution_unit_0_register_file_0_n_45_1));
	INV_X1_LVT execution_unit_0register_file_0i_45_2 (.A(execution_unit_0_register_file_0_n_45_1),.ZN(execution_unit_0_register_file_0_n_85));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_85),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_11 (.A1(execution_unit_0_register_file_0_r7[0]),.A2(execution_unit_0_register_file_0_n_83),.ZN(execution_unit_0_register_file_0_n_105_11));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_1 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r6_wr),.ZN(execution_unit_0_register_file_0_n_38_1));
	INV_X1_LVT execution_unit_0register_file_0i_38_2 (.A(execution_unit_0_register_file_0_n_38_1),.ZN(execution_unit_0_register_file_0_n_66));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_66),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_12 (.A1(execution_unit_0_register_file_0_r6[0]),.A2(execution_unit_0_register_file_0_n_64),.ZN(execution_unit_0_register_file_0_n_105_12));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_1 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r5_wr),.ZN(execution_unit_0_register_file_0_n_31_1));
	INV_X1_LVT execution_unit_0register_file_0i_31_2 (.A(execution_unit_0_register_file_0_n_31_1),.ZN(execution_unit_0_register_file_0_n_47));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_47),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_13 (.A1(execution_unit_0_register_file_0_r5[0]),.A2(execution_unit_0_register_file_0_n_45),.ZN(execution_unit_0_register_file_0_n_105_13));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_14 (.A1(execution_unit_0_register_file_0_n_105_10),.A2(execution_unit_0_register_file_0_n_105_11),.A3(execution_unit_0_register_file_0_n_105_12),.A4(execution_unit_0_register_file_0_n_105_13),.ZN(execution_unit_0_register_file_0_n_105_14));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_1 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r13_wr),.ZN(execution_unit_0_register_file_0_n_87_1));
	INV_X1_LVT execution_unit_0register_file_0i_87_2 (.A(execution_unit_0_register_file_0_n_87_1),.ZN(execution_unit_0_register_file_0_n_199));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_199),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[0]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_15 (.A1(execution_unit_0_register_file_0_r13[0]),.A2(execution_unit_0_register_file_0_n_197),.ZN(execution_unit_0_register_file_0_n_105_15));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_16 (.A1(execution_unit_0_register_file_0_n_105_4),.A2(execution_unit_0_register_file_0_n_105_9),.A3(execution_unit_0_register_file_0_n_105_14),.A4(execution_unit_0_register_file_0_n_105_15),.ZN(execution_unit_0_register_file_0_n_105_16));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_17 (.A1(pc[0]),.A2(execution_unit_0_register_file_0_n_254),.ZN(execution_unit_0_register_file_0_n_105_17));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_1 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r15_wr),.ZN(execution_unit_0_register_file_0_n_101_1));
	INV_X1_LVT execution_unit_0register_file_0i_101_2 (.A(execution_unit_0_register_file_0_n_101_1),.ZN(execution_unit_0_register_file_0_n_237));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_237),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_18 (.A1(execution_unit_0_register_file_0_r15[0]),.A2(execution_unit_0_register_file_0_n_235),.ZN(execution_unit_0_register_file_0_n_105_18));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_1 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[0]),.B1(execution_unit_0_alu_out[0]),.B2(execution_unit_0_register_file_0_r14_wr),.ZN(execution_unit_0_register_file_0_n_94_1));
	INV_X1_LVT execution_unit_0register_file_0i_94_2 (.A(execution_unit_0_register_file_0_n_94_1),.ZN(execution_unit_0_register_file_0_n_218));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b0___05F05d (.D(execution_unit_0_register_file_0_n_218),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[0]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_19 (.A1(execution_unit_0_register_file_0_r14[0]),.A2(execution_unit_0_register_file_0_n_216),.ZN(execution_unit_0_register_file_0_n_105_19));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_20 (.A1(execution_unit_0_register_file_0_n_105_16),.A2(execution_unit_0_register_file_0_n_105_17),.A3(execution_unit_0_register_file_0_n_105_18),.A4(execution_unit_0_register_file_0_n_105_19),.ZN(execution_unit_0_reg_src[0]));
	HA_X1_LVT execution_unit_0register_file_0i_22_0 (.A(execution_unit_0_register_file_0_n_25),.B(execution_unit_0_reg_src[0]),.CO(execution_unit_0_register_file_0_n_22_0),.S(execution_unit_0_register_file_0_reg_incr_val[0]));
	FA_X1_LVT execution_unit_0register_file_0i_22_1 (.A(execution_unit_0_register_file_0_n_26),.B(execution_unit_0_reg_src[1]),.CI(execution_unit_0_register_file_0_n_22_0),.CO(execution_unit_0_register_file_0_n_22_1),.S(execution_unit_0_register_file_0_reg_incr_val[1]));
	HA_X1_LVT execution_unit_0register_file_0i_22_2 (.A(execution_unit_0_reg_src[2]),.B(execution_unit_0_register_file_0_n_22_1),.CO(execution_unit_0_register_file_0_n_22_2),.S(execution_unit_0_register_file_0_reg_incr_val[2]));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_5 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_24_3));
	INV_X1_LVT execution_unit_0register_file_0i_24_6 (.A(execution_unit_0_register_file_0_n_24_3),.ZN(execution_unit_0_register_file_0_n_30));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_30),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_42 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[2]),.ZN(execution_unit_0_register_file_0_n_105_40));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b2___05F05d (.D(execution_unit_0_alu_out[2]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_43 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[2]),.ZN(execution_unit_0_register_file_0_n_105_41));
	INV_X1_LVT execution_unit_0register_file_0i_5_11 (.A(execution_unit_0_alu_stat_wr[2]),.ZN(execution_unit_0_register_file_0_n_5_9));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_12 (.A1(execution_unit_0_register_file_0_n_5_0),.A2(execution_unit_0_register_file_0_n_5_9),.A3(execution_unit_0_status[2]),.ZN(execution_unit_0_register_file_0_n_5_10));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_13 (.A1(execution_unit_0_register_file_0_n_5_9),.A2(execution_unit_0_register_file_0_r2_wr),.A3(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_5_11));
	NAND2_X1_LVT execution_unit_0register_file_0i_5_14 (.A1(execution_unit_0_alu_stat[2]),.A2(execution_unit_0_alu_stat_wr[2]),.ZN(execution_unit_0_register_file_0_n_5_12));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_15 (.A1(execution_unit_0_register_file_0_n_5_10),.A2(execution_unit_0_register_file_0_n_5_11),.A3(execution_unit_0_register_file_0_n_5_12),.ZN(execution_unit_0_register_file_0_n_11));
	AND2_X1_LVT execution_unit_0register_file_0i_6_3 (.A1(execution_unit_0_register_file_0_n_6_0),.A2(execution_unit_0_register_file_0_n_11),.ZN(execution_unit_0_register_file_0_n_15));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_15),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_status[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_44 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_status[2]),.ZN(execution_unit_0_register_file_0_n_105_42));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_2 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(execution_unit_0_alu_out[2]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[2]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_256),.ZN(execution_unit_0_register_file_0_n_109_1));
	INV_X1_LVT execution_unit_0register_file_0i_109_3 (.A(execution_unit_0_register_file_0_n_109_1),.ZN(execution_unit_0_register_file_0_n_274));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_274),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_45 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[2]),.ZN(execution_unit_0_register_file_0_n_105_43));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_46 (.A1(execution_unit_0_register_file_0_n_105_40),.A2(execution_unit_0_register_file_0_n_105_41),.A3(execution_unit_0_register_file_0_n_105_42),.A4(execution_unit_0_register_file_0_n_105_43),.ZN(execution_unit_0_register_file_0_n_105_44));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_5 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_80_3));
	INV_X1_LVT execution_unit_0register_file_0i_80_6 (.A(execution_unit_0_register_file_0_n_80_3),.ZN(execution_unit_0_register_file_0_n_182));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_182),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_47 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[2]),.ZN(execution_unit_0_register_file_0_n_105_45));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_5 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_73_3));
	INV_X1_LVT execution_unit_0register_file_0i_73_6 (.A(execution_unit_0_register_file_0_n_73_3),.ZN(execution_unit_0_register_file_0_n_163));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_163),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_48 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[2]),.ZN(execution_unit_0_register_file_0_n_105_46));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_5 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_66_3));
	INV_X1_LVT execution_unit_0register_file_0i_66_6 (.A(execution_unit_0_register_file_0_n_66_3),.ZN(execution_unit_0_register_file_0_n_144));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_144),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_49 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[2]),.ZN(execution_unit_0_register_file_0_n_105_47));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_5 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_59_3));
	INV_X1_LVT execution_unit_0register_file_0i_59_6 (.A(execution_unit_0_register_file_0_n_59_3),.ZN(execution_unit_0_register_file_0_n_125));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_125),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_50 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[2]),.ZN(execution_unit_0_register_file_0_n_105_48));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_51 (.A1(execution_unit_0_register_file_0_n_105_45),.A2(execution_unit_0_register_file_0_n_105_46),.A3(execution_unit_0_register_file_0_n_105_47),.A4(execution_unit_0_register_file_0_n_105_48),.ZN(execution_unit_0_register_file_0_n_105_49));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_5 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_52_3));
	INV_X1_LVT execution_unit_0register_file_0i_52_6 (.A(execution_unit_0_register_file_0_n_52_3),.ZN(execution_unit_0_register_file_0_n_106));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_106),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_52 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[2]),.ZN(execution_unit_0_register_file_0_n_105_50));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_5 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_45_3));
	INV_X1_LVT execution_unit_0register_file_0i_45_6 (.A(execution_unit_0_register_file_0_n_45_3),.ZN(execution_unit_0_register_file_0_n_87));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_87),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_53 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[2]),.ZN(execution_unit_0_register_file_0_n_105_51));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_5 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_38_3));
	INV_X1_LVT execution_unit_0register_file_0i_38_6 (.A(execution_unit_0_register_file_0_n_38_3),.ZN(execution_unit_0_register_file_0_n_68));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_68),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_54 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[2]),.ZN(execution_unit_0_register_file_0_n_105_52));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_5 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_31_3));
	INV_X1_LVT execution_unit_0register_file_0i_31_6 (.A(execution_unit_0_register_file_0_n_31_3),.ZN(execution_unit_0_register_file_0_n_49));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_49),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_55 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[2]),.ZN(execution_unit_0_register_file_0_n_105_53));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_56 (.A1(execution_unit_0_register_file_0_n_105_50),.A2(execution_unit_0_register_file_0_n_105_51),.A3(execution_unit_0_register_file_0_n_105_52),.A4(execution_unit_0_register_file_0_n_105_53),.ZN(execution_unit_0_register_file_0_n_105_54));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_5 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_87_3));
	INV_X1_LVT execution_unit_0register_file_0i_87_6 (.A(execution_unit_0_register_file_0_n_87_3),.ZN(execution_unit_0_register_file_0_n_201));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_201),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[2]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_57 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[2]),.ZN(execution_unit_0_register_file_0_n_105_55));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_58 (.A1(execution_unit_0_register_file_0_n_105_44),.A2(execution_unit_0_register_file_0_n_105_49),.A3(execution_unit_0_register_file_0_n_105_54),.A4(execution_unit_0_register_file_0_n_105_55),.ZN(execution_unit_0_register_file_0_n_105_56));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_59 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[2]),.ZN(execution_unit_0_register_file_0_n_105_57));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_5 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_101_3));
	INV_X1_LVT execution_unit_0register_file_0i_101_6 (.A(execution_unit_0_register_file_0_n_101_3),.ZN(execution_unit_0_register_file_0_n_239));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_239),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_60 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[2]),.ZN(execution_unit_0_register_file_0_n_105_58));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_5 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[2]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(execution_unit_0_alu_out[2]),.ZN(execution_unit_0_register_file_0_n_94_3));
	INV_X1_LVT execution_unit_0register_file_0i_94_6 (.A(execution_unit_0_register_file_0_n_94_3),.ZN(execution_unit_0_register_file_0_n_220));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b2___05F05d (.D(execution_unit_0_register_file_0_n_220),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[2]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_61 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[2]),.ZN(execution_unit_0_register_file_0_n_105_59));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_62 (.A1(execution_unit_0_register_file_0_n_105_56),.A2(execution_unit_0_register_file_0_n_105_57),.A3(execution_unit_0_register_file_0_n_105_58),.A4(execution_unit_0_register_file_0_n_105_59),.ZN(execution_unit_0_reg_src[2]));
	HA_X1_LVT execution_unit_0register_file_0i_106_1 (.A(execution_unit_0_reg_src[2]),.B(execution_unit_0_reg_src[1]),.CO(execution_unit_0_register_file_0_n_106_0),.S(execution_unit_0_register_file_0_n_256));
	HA_X1_LVT execution_unit_0register_file_0i_106_2 (.A(execution_unit_0_reg_src[3]),.B(execution_unit_0_register_file_0_n_106_0),.CO(execution_unit_0_register_file_0_n_106_1),.S(execution_unit_0_register_file_0_n_257));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_4 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(execution_unit_0_alu_out[3]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[3]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_257),.ZN(execution_unit_0_register_file_0_n_109_2));
	INV_X1_LVT execution_unit_0register_file_0i_109_5 (.A(execution_unit_0_register_file_0_n_109_2),.ZN(execution_unit_0_register_file_0_n_275));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_275),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_66 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[3]),.ZN(execution_unit_0_register_file_0_n_105_63));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_67 (.A1(execution_unit_0_register_file_0_n_105_60),.A2(execution_unit_0_register_file_0_n_105_61),.A3(execution_unit_0_register_file_0_n_105_62),.A4(execution_unit_0_register_file_0_n_105_63),.ZN(execution_unit_0_register_file_0_n_105_64));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_7 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_80_4));
	INV_X1_LVT execution_unit_0register_file_0i_80_8 (.A(execution_unit_0_register_file_0_n_80_4),.ZN(execution_unit_0_register_file_0_n_183));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_183),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_68 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[3]),.ZN(execution_unit_0_register_file_0_n_105_65));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_7 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_73_4));
	INV_X1_LVT execution_unit_0register_file_0i_73_8 (.A(execution_unit_0_register_file_0_n_73_4),.ZN(execution_unit_0_register_file_0_n_164));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_164),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_69 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[3]),.ZN(execution_unit_0_register_file_0_n_105_66));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_7 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_66_4));
	INV_X1_LVT execution_unit_0register_file_0i_66_8 (.A(execution_unit_0_register_file_0_n_66_4),.ZN(execution_unit_0_register_file_0_n_145));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_145),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_70 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[3]),.ZN(execution_unit_0_register_file_0_n_105_67));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_7 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_59_4));
	INV_X1_LVT execution_unit_0register_file_0i_59_8 (.A(execution_unit_0_register_file_0_n_59_4),.ZN(execution_unit_0_register_file_0_n_126));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_126),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_71 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[3]),.ZN(execution_unit_0_register_file_0_n_105_68));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_72 (.A1(execution_unit_0_register_file_0_n_105_65),.A2(execution_unit_0_register_file_0_n_105_66),.A3(execution_unit_0_register_file_0_n_105_67),.A4(execution_unit_0_register_file_0_n_105_68),.ZN(execution_unit_0_register_file_0_n_105_69));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_7 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_52_4));
	INV_X1_LVT execution_unit_0register_file_0i_52_8 (.A(execution_unit_0_register_file_0_n_52_4),.ZN(execution_unit_0_register_file_0_n_107));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_107),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_73 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[3]),.ZN(execution_unit_0_register_file_0_n_105_70));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_7 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_45_4));
	INV_X1_LVT execution_unit_0register_file_0i_45_8 (.A(execution_unit_0_register_file_0_n_45_4),.ZN(execution_unit_0_register_file_0_n_88));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_88),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_74 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[3]),.ZN(execution_unit_0_register_file_0_n_105_71));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_7 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_38_4));
	INV_X1_LVT execution_unit_0register_file_0i_38_8 (.A(execution_unit_0_register_file_0_n_38_4),.ZN(execution_unit_0_register_file_0_n_69));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_69),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_75 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[3]),.ZN(execution_unit_0_register_file_0_n_105_72));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_7 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_31_4));
	INV_X1_LVT execution_unit_0register_file_0i_31_8 (.A(execution_unit_0_register_file_0_n_31_4),.ZN(execution_unit_0_register_file_0_n_50));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_50),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_76 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[3]),.ZN(execution_unit_0_register_file_0_n_105_73));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_77 (.A1(execution_unit_0_register_file_0_n_105_70),.A2(execution_unit_0_register_file_0_n_105_71),.A3(execution_unit_0_register_file_0_n_105_72),.A4(execution_unit_0_register_file_0_n_105_73),.ZN(execution_unit_0_register_file_0_n_105_74));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_7 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_87_4));
	INV_X1_LVT execution_unit_0register_file_0i_87_8 (.A(execution_unit_0_register_file_0_n_87_4),.ZN(execution_unit_0_register_file_0_n_202));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_202),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[3]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_78 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[3]),.ZN(execution_unit_0_register_file_0_n_105_75));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_79 (.A1(execution_unit_0_register_file_0_n_105_64),.A2(execution_unit_0_register_file_0_n_105_69),.A3(execution_unit_0_register_file_0_n_105_74),.A4(execution_unit_0_register_file_0_n_105_75),.ZN(execution_unit_0_register_file_0_n_105_76));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_80 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[3]),.ZN(execution_unit_0_register_file_0_n_105_77));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_7 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_101_4));
	INV_X1_LVT execution_unit_0register_file_0i_101_8 (.A(execution_unit_0_register_file_0_n_101_4),.ZN(execution_unit_0_register_file_0_n_240));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_240),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_81 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[3]),.ZN(execution_unit_0_register_file_0_n_105_78));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_7 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[3]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(execution_unit_0_alu_out[3]),.ZN(execution_unit_0_register_file_0_n_94_4));
	INV_X1_LVT execution_unit_0register_file_0i_94_8 (.A(execution_unit_0_register_file_0_n_94_4),.ZN(execution_unit_0_register_file_0_n_221));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b3___05F05d (.D(execution_unit_0_register_file_0_n_221),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_82 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[3]),.ZN(execution_unit_0_register_file_0_n_105_79));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_83 (.A1(execution_unit_0_register_file_0_n_105_76),.A2(execution_unit_0_register_file_0_n_105_77),.A3(execution_unit_0_register_file_0_n_105_78),.A4(execution_unit_0_register_file_0_n_105_79),.ZN(execution_unit_0_reg_src[3]));
	HA_X1_LVT execution_unit_0register_file_0i_22_3 (.A(execution_unit_0_reg_src[3]),.B(execution_unit_0_register_file_0_n_22_2),.CO(execution_unit_0_register_file_0_n_22_3),.S(execution_unit_0_register_file_0_reg_incr_val[3]));
	HA_X1_LVT execution_unit_0register_file_0i_22_4 (.A(execution_unit_0_reg_src[4]),.B(execution_unit_0_register_file_0_n_22_3),.CO(execution_unit_0_register_file_0_n_22_4),.S(execution_unit_0_register_file_0_reg_incr_val[4]));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_9 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_24_5));
	INV_X1_LVT execution_unit_0register_file_0i_24_10 (.A(execution_unit_0_register_file_0_n_24_5),.ZN(execution_unit_0_register_file_0_n_32));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_32),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_84 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[4]),.ZN(execution_unit_0_register_file_0_n_105_80));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b4___05F05d (.D(execution_unit_0_alu_out[4]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_85 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[4]),.ZN(execution_unit_0_register_file_0_n_105_81));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_86 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_register_file_0_n_7),.ZN(execution_unit_0_register_file_0_n_105_82));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_6 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(execution_unit_0_alu_out[4]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[4]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_258),.ZN(execution_unit_0_register_file_0_n_109_3));
	INV_X1_LVT execution_unit_0register_file_0i_109_7 (.A(execution_unit_0_register_file_0_n_109_3),.ZN(execution_unit_0_register_file_0_n_276));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_276),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_87 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[4]),.ZN(execution_unit_0_register_file_0_n_105_83));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_88 (.A1(execution_unit_0_register_file_0_n_105_80),.A2(execution_unit_0_register_file_0_n_105_81),.A3(execution_unit_0_register_file_0_n_105_82),.A4(execution_unit_0_register_file_0_n_105_83),.ZN(execution_unit_0_register_file_0_n_105_84));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_9 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_80_5));
	INV_X1_LVT execution_unit_0register_file_0i_80_10 (.A(execution_unit_0_register_file_0_n_80_5),.ZN(execution_unit_0_register_file_0_n_184));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_184),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_89 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[4]),.ZN(execution_unit_0_register_file_0_n_105_85));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_9 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_73_5));
	INV_X1_LVT execution_unit_0register_file_0i_73_10 (.A(execution_unit_0_register_file_0_n_73_5),.ZN(execution_unit_0_register_file_0_n_165));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_165),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_90 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[4]),.ZN(execution_unit_0_register_file_0_n_105_86));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_9 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_66_5));
	INV_X1_LVT execution_unit_0register_file_0i_66_10 (.A(execution_unit_0_register_file_0_n_66_5),.ZN(execution_unit_0_register_file_0_n_146));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_146),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_91 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[4]),.ZN(execution_unit_0_register_file_0_n_105_87));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_9 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_59_5));
	INV_X1_LVT execution_unit_0register_file_0i_59_10 (.A(execution_unit_0_register_file_0_n_59_5),.ZN(execution_unit_0_register_file_0_n_127));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_127),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_92 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[4]),.ZN(execution_unit_0_register_file_0_n_105_88));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_93 (.A1(execution_unit_0_register_file_0_n_105_85),.A2(execution_unit_0_register_file_0_n_105_86),.A3(execution_unit_0_register_file_0_n_105_87),.A4(execution_unit_0_register_file_0_n_105_88),.ZN(execution_unit_0_register_file_0_n_105_89));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_9 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_52_5));
	INV_X1_LVT execution_unit_0register_file_0i_52_10 (.A(execution_unit_0_register_file_0_n_52_5),.ZN(execution_unit_0_register_file_0_n_108));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_108),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_94 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[4]),.ZN(execution_unit_0_register_file_0_n_105_90));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_9 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_45_5));
	INV_X1_LVT execution_unit_0register_file_0i_45_10 (.A(execution_unit_0_register_file_0_n_45_5),.ZN(execution_unit_0_register_file_0_n_89));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_89),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_95 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[4]),.ZN(execution_unit_0_register_file_0_n_105_91));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_9 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_38_5));
	INV_X1_LVT execution_unit_0register_file_0i_38_10 (.A(execution_unit_0_register_file_0_n_38_5),.ZN(execution_unit_0_register_file_0_n_70));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_70),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_96 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[4]),.ZN(execution_unit_0_register_file_0_n_105_92));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_9 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_31_5));
	INV_X1_LVT execution_unit_0register_file_0i_31_10 (.A(execution_unit_0_register_file_0_n_31_5),.ZN(execution_unit_0_register_file_0_n_51));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_51),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_97 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[4]),.ZN(execution_unit_0_register_file_0_n_105_93));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_98 (.A1(execution_unit_0_register_file_0_n_105_90),.A2(execution_unit_0_register_file_0_n_105_91),.A3(execution_unit_0_register_file_0_n_105_92),.A4(execution_unit_0_register_file_0_n_105_93),.ZN(execution_unit_0_register_file_0_n_105_94));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_9 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_87_5));
	INV_X1_LVT execution_unit_0register_file_0i_87_10 (.A(execution_unit_0_register_file_0_n_87_5),.ZN(execution_unit_0_register_file_0_n_203));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_203),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[4]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_99 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[4]),.ZN(execution_unit_0_register_file_0_n_105_95));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_100 (.A1(execution_unit_0_register_file_0_n_105_84),.A2(execution_unit_0_register_file_0_n_105_89),.A3(execution_unit_0_register_file_0_n_105_94),.A4(execution_unit_0_register_file_0_n_105_95),.ZN(execution_unit_0_register_file_0_n_105_96));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_101 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[4]),.ZN(execution_unit_0_register_file_0_n_105_97));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_9 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_101_5));
	INV_X1_LVT execution_unit_0register_file_0i_101_10 (.A(execution_unit_0_register_file_0_n_101_5),.ZN(execution_unit_0_register_file_0_n_241));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_241),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_102 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[4]),.ZN(execution_unit_0_register_file_0_n_105_98));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_9 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[4]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(execution_unit_0_alu_out[4]),.ZN(execution_unit_0_register_file_0_n_94_5));
	INV_X1_LVT execution_unit_0register_file_0i_94_10 (.A(execution_unit_0_register_file_0_n_94_5),.ZN(execution_unit_0_register_file_0_n_222));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b4___05F05d (.D(execution_unit_0_register_file_0_n_222),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[4]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_103 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[4]),.ZN(execution_unit_0_register_file_0_n_105_99));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_104 (.A1(execution_unit_0_register_file_0_n_105_96),.A2(execution_unit_0_register_file_0_n_105_97),.A3(execution_unit_0_register_file_0_n_105_98),.A4(execution_unit_0_register_file_0_n_105_99),.ZN(execution_unit_0_reg_src[4]));
	HA_X1_LVT execution_unit_0register_file_0i_106_3 (.A(execution_unit_0_reg_src[4]),.B(execution_unit_0_register_file_0_n_106_1),.CO(execution_unit_0_register_file_0_n_106_2),.S(execution_unit_0_register_file_0_n_258));
	HA_X1_LVT execution_unit_0register_file_0i_106_4 (.A(execution_unit_0_reg_src[5]),.B(execution_unit_0_register_file_0_n_106_2),.CO(execution_unit_0_register_file_0_n_106_3),.S(execution_unit_0_register_file_0_n_259));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_8 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(execution_unit_0_alu_out[5]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[5]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_259),.ZN(execution_unit_0_register_file_0_n_109_4));
	INV_X1_LVT execution_unit_0register_file_0i_109_9 (.A(execution_unit_0_register_file_0_n_109_4),.ZN(execution_unit_0_register_file_0_n_277));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_277),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_108 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[5]),.ZN(execution_unit_0_register_file_0_n_105_103));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_109 (.A1(execution_unit_0_register_file_0_n_105_100),.A2(execution_unit_0_register_file_0_n_105_101),.A3(execution_unit_0_register_file_0_n_105_102),.A4(execution_unit_0_register_file_0_n_105_103),.ZN(execution_unit_0_register_file_0_n_105_104));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_11 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_80_6));
	INV_X1_LVT execution_unit_0register_file_0i_80_12 (.A(execution_unit_0_register_file_0_n_80_6),.ZN(execution_unit_0_register_file_0_n_185));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_185),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_110 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[5]),.ZN(execution_unit_0_register_file_0_n_105_105));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_11 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_73_6));
	INV_X1_LVT execution_unit_0register_file_0i_73_12 (.A(execution_unit_0_register_file_0_n_73_6),.ZN(execution_unit_0_register_file_0_n_166));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_166),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_111 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[5]),.ZN(execution_unit_0_register_file_0_n_105_106));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_11 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_66_6));
	INV_X1_LVT execution_unit_0register_file_0i_66_12 (.A(execution_unit_0_register_file_0_n_66_6),.ZN(execution_unit_0_register_file_0_n_147));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_147),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_112 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[5]),.ZN(execution_unit_0_register_file_0_n_105_107));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_11 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_59_6));
	INV_X1_LVT execution_unit_0register_file_0i_59_12 (.A(execution_unit_0_register_file_0_n_59_6),.ZN(execution_unit_0_register_file_0_n_128));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_128),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_113 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[5]),.ZN(execution_unit_0_register_file_0_n_105_108));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_114 (.A1(execution_unit_0_register_file_0_n_105_105),.A2(execution_unit_0_register_file_0_n_105_106),.A3(execution_unit_0_register_file_0_n_105_107),.A4(execution_unit_0_register_file_0_n_105_108),.ZN(execution_unit_0_register_file_0_n_105_109));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_11 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_52_6));
	INV_X1_LVT execution_unit_0register_file_0i_52_12 (.A(execution_unit_0_register_file_0_n_52_6),.ZN(execution_unit_0_register_file_0_n_109));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_109),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_115 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[5]),.ZN(execution_unit_0_register_file_0_n_105_110));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_11 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_45_6));
	INV_X1_LVT execution_unit_0register_file_0i_45_12 (.A(execution_unit_0_register_file_0_n_45_6),.ZN(execution_unit_0_register_file_0_n_90));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_90),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_116 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[5]),.ZN(execution_unit_0_register_file_0_n_105_111));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_11 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_38_6));
	INV_X1_LVT execution_unit_0register_file_0i_38_12 (.A(execution_unit_0_register_file_0_n_38_6),.ZN(execution_unit_0_register_file_0_n_71));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_71),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_117 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[5]),.ZN(execution_unit_0_register_file_0_n_105_112));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_11 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_31_6));
	INV_X1_LVT execution_unit_0register_file_0i_31_12 (.A(execution_unit_0_register_file_0_n_31_6),.ZN(execution_unit_0_register_file_0_n_52));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_52),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_118 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[5]),.ZN(execution_unit_0_register_file_0_n_105_113));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_119 (.A1(execution_unit_0_register_file_0_n_105_110),.A2(execution_unit_0_register_file_0_n_105_111),.A3(execution_unit_0_register_file_0_n_105_112),.A4(execution_unit_0_register_file_0_n_105_113),.ZN(execution_unit_0_register_file_0_n_105_114));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_11 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_87_6));
	INV_X1_LVT execution_unit_0register_file_0i_87_12 (.A(execution_unit_0_register_file_0_n_87_6),.ZN(execution_unit_0_register_file_0_n_204));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_204),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[5]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_120 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[5]),.ZN(execution_unit_0_register_file_0_n_105_115));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_121 (.A1(execution_unit_0_register_file_0_n_105_104),.A2(execution_unit_0_register_file_0_n_105_109),.A3(execution_unit_0_register_file_0_n_105_114),.A4(execution_unit_0_register_file_0_n_105_115),.ZN(execution_unit_0_register_file_0_n_105_116));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_122 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[5]),.ZN(execution_unit_0_register_file_0_n_105_117));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_11 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_101_6));
	INV_X1_LVT execution_unit_0register_file_0i_101_12 (.A(execution_unit_0_register_file_0_n_101_6),.ZN(execution_unit_0_register_file_0_n_242));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_242),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_123 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[5]),.ZN(execution_unit_0_register_file_0_n_105_118));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_11 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[5]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(execution_unit_0_alu_out[5]),.ZN(execution_unit_0_register_file_0_n_94_6));
	INV_X1_LVT execution_unit_0register_file_0i_94_12 (.A(execution_unit_0_register_file_0_n_94_6),.ZN(execution_unit_0_register_file_0_n_223));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b5___05F05d (.D(execution_unit_0_register_file_0_n_223),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[5]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_124 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[5]),.ZN(execution_unit_0_register_file_0_n_105_119));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_125 (.A1(execution_unit_0_register_file_0_n_105_116),.A2(execution_unit_0_register_file_0_n_105_117),.A3(execution_unit_0_register_file_0_n_105_118),.A4(execution_unit_0_register_file_0_n_105_119),.ZN(execution_unit_0_reg_src[5]));
	HA_X1_LVT execution_unit_0register_file_0i_22_5 (.A(execution_unit_0_reg_src[5]),.B(execution_unit_0_register_file_0_n_22_4),.CO(execution_unit_0_register_file_0_n_22_5),.S(execution_unit_0_register_file_0_reg_incr_val[5]));
	HA_X1_LVT execution_unit_0register_file_0i_22_6 (.A(execution_unit_0_reg_src[6]),.B(execution_unit_0_register_file_0_n_22_5),.CO(execution_unit_0_register_file_0_n_22_6),.S(execution_unit_0_register_file_0_reg_incr_val[6]));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_13 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_24_7));
	INV_X1_LVT execution_unit_0register_file_0i_24_14 (.A(execution_unit_0_register_file_0_n_24_7),.ZN(execution_unit_0_register_file_0_n_34));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_34),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_126 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[6]),.ZN(execution_unit_0_register_file_0_n_105_120));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b6___05F05d (.D(execution_unit_0_alu_out[6]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_127 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[6]),.ZN(execution_unit_0_register_file_0_n_105_121));
	AOI22_X1_LVT execution_unit_0register_file_0i_2_5 (.A1(execution_unit_0_register_file_0_n_2_0),.A2(scg0),.B1(execution_unit_0_register_file_0_r2_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_2_3));
	INV_X1_LVT execution_unit_0register_file_0i_2_6 (.A(execution_unit_0_register_file_0_n_2_3),.ZN(execution_unit_0_register_file_0_r2_nxt[3]));
	AND2_X1_LVT execution_unit_0register_file_0i_6_6 (.A1(execution_unit_0_register_file_0_n_6_0),.A2(execution_unit_0_register_file_0_r2_nxt[3]),.ZN(execution_unit_0_register_file_0_n_18));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_18),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(scg0),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_128 (.A1(execution_unit_0_register_file_0_n_21),.A2(scg0),.ZN(execution_unit_0_register_file_0_n_105_122));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_10 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(execution_unit_0_alu_out[6]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[6]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_260),.ZN(execution_unit_0_register_file_0_n_109_5));
	INV_X1_LVT execution_unit_0register_file_0i_109_11 (.A(execution_unit_0_register_file_0_n_109_5),.ZN(execution_unit_0_register_file_0_n_278));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_278),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_129 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[6]),.ZN(execution_unit_0_register_file_0_n_105_123));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_130 (.A1(execution_unit_0_register_file_0_n_105_120),.A2(execution_unit_0_register_file_0_n_105_121),.A3(execution_unit_0_register_file_0_n_105_122),.A4(execution_unit_0_register_file_0_n_105_123),.ZN(execution_unit_0_register_file_0_n_105_124));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_13 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_80_7));
	INV_X1_LVT execution_unit_0register_file_0i_80_14 (.A(execution_unit_0_register_file_0_n_80_7),.ZN(execution_unit_0_register_file_0_n_186));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_186),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_131 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[6]),.ZN(execution_unit_0_register_file_0_n_105_125));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_13 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_73_7));
	INV_X1_LVT execution_unit_0register_file_0i_73_14 (.A(execution_unit_0_register_file_0_n_73_7),.ZN(execution_unit_0_register_file_0_n_167));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_167),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_132 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[6]),.ZN(execution_unit_0_register_file_0_n_105_126));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_13 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_66_7));
	INV_X1_LVT execution_unit_0register_file_0i_66_14 (.A(execution_unit_0_register_file_0_n_66_7),.ZN(execution_unit_0_register_file_0_n_148));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_148),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_133 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[6]),.ZN(execution_unit_0_register_file_0_n_105_127));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_13 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_59_7));
	INV_X1_LVT execution_unit_0register_file_0i_59_14 (.A(execution_unit_0_register_file_0_n_59_7),.ZN(execution_unit_0_register_file_0_n_129));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_129),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_134 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[6]),.ZN(execution_unit_0_register_file_0_n_105_128));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_135 (.A1(execution_unit_0_register_file_0_n_105_125),.A2(execution_unit_0_register_file_0_n_105_126),.A3(execution_unit_0_register_file_0_n_105_127),.A4(execution_unit_0_register_file_0_n_105_128),.ZN(execution_unit_0_register_file_0_n_105_129));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_13 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_52_7));
	INV_X1_LVT execution_unit_0register_file_0i_52_14 (.A(execution_unit_0_register_file_0_n_52_7),.ZN(execution_unit_0_register_file_0_n_110));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_110),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_136 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[6]),.ZN(execution_unit_0_register_file_0_n_105_130));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_13 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_45_7));
	INV_X1_LVT execution_unit_0register_file_0i_45_14 (.A(execution_unit_0_register_file_0_n_45_7),.ZN(execution_unit_0_register_file_0_n_91));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_91),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_137 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[6]),.ZN(execution_unit_0_register_file_0_n_105_131));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_13 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_38_7));
	INV_X1_LVT execution_unit_0register_file_0i_38_14 (.A(execution_unit_0_register_file_0_n_38_7),.ZN(execution_unit_0_register_file_0_n_72));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_72),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_138 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[6]),.ZN(execution_unit_0_register_file_0_n_105_132));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_13 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_31_7));
	INV_X1_LVT execution_unit_0register_file_0i_31_14 (.A(execution_unit_0_register_file_0_n_31_7),.ZN(execution_unit_0_register_file_0_n_53));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_53),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_139 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[6]),.ZN(execution_unit_0_register_file_0_n_105_133));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_140 (.A1(execution_unit_0_register_file_0_n_105_130),.A2(execution_unit_0_register_file_0_n_105_131),.A3(execution_unit_0_register_file_0_n_105_132),.A4(execution_unit_0_register_file_0_n_105_133),.ZN(execution_unit_0_register_file_0_n_105_134));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_13 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_87_7));
	INV_X1_LVT execution_unit_0register_file_0i_87_14 (.A(execution_unit_0_register_file_0_n_87_7),.ZN(execution_unit_0_register_file_0_n_205));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_205),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[6]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_141 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[6]),.ZN(execution_unit_0_register_file_0_n_105_135));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_142 (.A1(execution_unit_0_register_file_0_n_105_124),.A2(execution_unit_0_register_file_0_n_105_129),.A3(execution_unit_0_register_file_0_n_105_134),.A4(execution_unit_0_register_file_0_n_105_135),.ZN(execution_unit_0_register_file_0_n_105_136));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_143 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[6]),.ZN(execution_unit_0_register_file_0_n_105_137));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_13 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_101_7));
	INV_X1_LVT execution_unit_0register_file_0i_101_14 (.A(execution_unit_0_register_file_0_n_101_7),.ZN(execution_unit_0_register_file_0_n_243));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_243),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_144 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[6]),.ZN(execution_unit_0_register_file_0_n_105_138));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_13 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[6]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(execution_unit_0_alu_out[6]),.ZN(execution_unit_0_register_file_0_n_94_7));
	INV_X1_LVT execution_unit_0register_file_0i_94_14 (.A(execution_unit_0_register_file_0_n_94_7),.ZN(execution_unit_0_register_file_0_n_224));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b6___05F05d (.D(execution_unit_0_register_file_0_n_224),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[6]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_145 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[6]),.ZN(execution_unit_0_register_file_0_n_105_139));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_146 (.A1(execution_unit_0_register_file_0_n_105_136),.A2(execution_unit_0_register_file_0_n_105_137),.A3(execution_unit_0_register_file_0_n_105_138),.A4(execution_unit_0_register_file_0_n_105_139),.ZN(execution_unit_0_reg_src[6]));
	HA_X1_LVT execution_unit_0register_file_0i_106_5 (.A(execution_unit_0_reg_src[6]),.B(execution_unit_0_register_file_0_n_106_3),.CO(execution_unit_0_register_file_0_n_106_4),.S(execution_unit_0_register_file_0_n_260));
	HA_X1_LVT execution_unit_0register_file_0i_106_6 (.A(execution_unit_0_reg_src[7]),.B(execution_unit_0_register_file_0_n_106_4),.CO(execution_unit_0_register_file_0_n_106_5),.S(execution_unit_0_register_file_0_n_261));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_12 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(execution_unit_0_alu_out[7]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[7]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_261),.ZN(execution_unit_0_register_file_0_n_109_6));
	INV_X1_LVT execution_unit_0register_file_0i_109_13 (.A(execution_unit_0_register_file_0_n_109_6),.ZN(execution_unit_0_register_file_0_n_279));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_279),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_150 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[7]),.ZN(execution_unit_0_register_file_0_n_105_143));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_151 (.A1(execution_unit_0_register_file_0_n_105_140),.A2(execution_unit_0_register_file_0_n_105_141),.A3(execution_unit_0_register_file_0_n_105_142),.A4(execution_unit_0_register_file_0_n_105_143),.ZN(execution_unit_0_register_file_0_n_105_144));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_15 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_80_8));
	INV_X1_LVT execution_unit_0register_file_0i_80_16 (.A(execution_unit_0_register_file_0_n_80_8),.ZN(execution_unit_0_register_file_0_n_187));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_187),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_152 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[7]),.ZN(execution_unit_0_register_file_0_n_105_145));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_15 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_73_8));
	INV_X1_LVT execution_unit_0register_file_0i_73_16 (.A(execution_unit_0_register_file_0_n_73_8),.ZN(execution_unit_0_register_file_0_n_168));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_168),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_153 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[7]),.ZN(execution_unit_0_register_file_0_n_105_146));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_15 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_66_8));
	INV_X1_LVT execution_unit_0register_file_0i_66_16 (.A(execution_unit_0_register_file_0_n_66_8),.ZN(execution_unit_0_register_file_0_n_149));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_149),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_154 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[7]),.ZN(execution_unit_0_register_file_0_n_105_147));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_15 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_59_8));
	INV_X1_LVT execution_unit_0register_file_0i_59_16 (.A(execution_unit_0_register_file_0_n_59_8),.ZN(execution_unit_0_register_file_0_n_130));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_130),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_155 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[7]),.ZN(execution_unit_0_register_file_0_n_105_148));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_156 (.A1(execution_unit_0_register_file_0_n_105_145),.A2(execution_unit_0_register_file_0_n_105_146),.A3(execution_unit_0_register_file_0_n_105_147),.A4(execution_unit_0_register_file_0_n_105_148),.ZN(execution_unit_0_register_file_0_n_105_149));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_15 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_52_8));
	INV_X1_LVT execution_unit_0register_file_0i_52_16 (.A(execution_unit_0_register_file_0_n_52_8),.ZN(execution_unit_0_register_file_0_n_111));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_111),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_157 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[7]),.ZN(execution_unit_0_register_file_0_n_105_150));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_15 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_45_8));
	INV_X1_LVT execution_unit_0register_file_0i_45_16 (.A(execution_unit_0_register_file_0_n_45_8),.ZN(execution_unit_0_register_file_0_n_92));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_92),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_158 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[7]),.ZN(execution_unit_0_register_file_0_n_105_151));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_15 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_38_8));
	INV_X1_LVT execution_unit_0register_file_0i_38_16 (.A(execution_unit_0_register_file_0_n_38_8),.ZN(execution_unit_0_register_file_0_n_73));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_73),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_159 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[7]),.ZN(execution_unit_0_register_file_0_n_105_152));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_15 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_31_8));
	INV_X1_LVT execution_unit_0register_file_0i_31_16 (.A(execution_unit_0_register_file_0_n_31_8),.ZN(execution_unit_0_register_file_0_n_54));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_54),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_160 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[7]),.ZN(execution_unit_0_register_file_0_n_105_153));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_161 (.A1(execution_unit_0_register_file_0_n_105_150),.A2(execution_unit_0_register_file_0_n_105_151),.A3(execution_unit_0_register_file_0_n_105_152),.A4(execution_unit_0_register_file_0_n_105_153),.ZN(execution_unit_0_register_file_0_n_105_154));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_15 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_87_8));
	INV_X1_LVT execution_unit_0register_file_0i_87_16 (.A(execution_unit_0_register_file_0_n_87_8),.ZN(execution_unit_0_register_file_0_n_206));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_206),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[7]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_162 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[7]),.ZN(execution_unit_0_register_file_0_n_105_155));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_163 (.A1(execution_unit_0_register_file_0_n_105_144),.A2(execution_unit_0_register_file_0_n_105_149),.A3(execution_unit_0_register_file_0_n_105_154),.A4(execution_unit_0_register_file_0_n_105_155),.ZN(execution_unit_0_register_file_0_n_105_156));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_164 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[7]),.ZN(execution_unit_0_register_file_0_n_105_157));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_15 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_101_8));
	INV_X1_LVT execution_unit_0register_file_0i_101_16 (.A(execution_unit_0_register_file_0_n_101_8),.ZN(execution_unit_0_register_file_0_n_244));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_244),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_165 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[7]),.ZN(execution_unit_0_register_file_0_n_105_158));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_15 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[7]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(execution_unit_0_alu_out[7]),.ZN(execution_unit_0_register_file_0_n_94_8));
	INV_X1_LVT execution_unit_0register_file_0i_94_16 (.A(execution_unit_0_register_file_0_n_94_8),.ZN(execution_unit_0_register_file_0_n_225));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b7___05F05d (.D(execution_unit_0_register_file_0_n_225),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[7]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_166 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[7]),.ZN(execution_unit_0_register_file_0_n_105_159));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_167 (.A1(execution_unit_0_register_file_0_n_105_156),.A2(execution_unit_0_register_file_0_n_105_157),.A3(execution_unit_0_register_file_0_n_105_158),.A4(execution_unit_0_register_file_0_n_105_159),.ZN(execution_unit_0_reg_src[7]));
	HA_X1_LVT execution_unit_0register_file_0i_22_7 (.A(execution_unit_0_reg_src[7]),.B(execution_unit_0_register_file_0_n_22_6),.CO(execution_unit_0_register_file_0_n_22_7),.S(execution_unit_0_register_file_0_reg_incr_val[7]));
	HA_X1_LVT execution_unit_0register_file_0i_22_8 (.A(execution_unit_0_reg_src[8]),.B(execution_unit_0_register_file_0_n_22_7),.CO(execution_unit_0_register_file_0_n_22_8),.S(execution_unit_0_register_file_0_reg_incr_val[8]));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_17 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_24_9));
	INV_X1_LVT execution_unit_0register_file_0i_24_18 (.A(execution_unit_0_register_file_0_n_24_9),.ZN(execution_unit_0_register_file_0_n_36));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_36),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_168 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[8]),.ZN(execution_unit_0_register_file_0_n_105_160));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b8___05F05d (.D(pc_sw[8]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_169 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[8]),.ZN(execution_unit_0_register_file_0_n_105_161));
	INV_X1_LVT execution_unit_0register_file_0i_5_16 (.A(execution_unit_0_alu_stat_wr[3]),.ZN(execution_unit_0_register_file_0_n_5_13));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_17 (.A1(execution_unit_0_register_file_0_n_5_0),.A2(execution_unit_0_register_file_0_n_5_13),.A3(execution_unit_0_status[3]),.ZN(execution_unit_0_register_file_0_n_5_14));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_18 (.A1(execution_unit_0_register_file_0_n_5_13),.A2(execution_unit_0_register_file_0_r2_wr),.A3(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_5_15));
	NAND2_X1_LVT execution_unit_0register_file_0i_5_19 (.A1(execution_unit_0_alu_stat[3]),.A2(execution_unit_0_alu_stat_wr[3]),.ZN(execution_unit_0_register_file_0_n_5_16));
	NAND3_X1_LVT execution_unit_0register_file_0i_5_20 (.A1(execution_unit_0_register_file_0_n_5_14),.A2(execution_unit_0_register_file_0_n_5_15),.A3(execution_unit_0_register_file_0_n_5_16),.ZN(execution_unit_0_register_file_0_n_12));
	AND2_X1_LVT execution_unit_0register_file_0i_6_8 (.A1(execution_unit_0_register_file_0_n_6_0),.A2(execution_unit_0_register_file_0_n_12),.ZN(execution_unit_0_register_file_0_n_20));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_20),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_status[3]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_170 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_status[3]),.ZN(execution_unit_0_register_file_0_n_105_162));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_14 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(pc_sw[8]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[8]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_262),.ZN(execution_unit_0_register_file_0_n_109_7));
	INV_X1_LVT execution_unit_0register_file_0i_109_15 (.A(execution_unit_0_register_file_0_n_109_7),.ZN(execution_unit_0_register_file_0_n_280));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_280),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_171 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[8]),.ZN(execution_unit_0_register_file_0_n_105_163));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_172 (.A1(execution_unit_0_register_file_0_n_105_160),.A2(execution_unit_0_register_file_0_n_105_161),.A3(execution_unit_0_register_file_0_n_105_162),.A4(execution_unit_0_register_file_0_n_105_163),.ZN(execution_unit_0_register_file_0_n_105_164));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_17 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_80_9));
	INV_X1_LVT execution_unit_0register_file_0i_80_18 (.A(execution_unit_0_register_file_0_n_80_9),.ZN(execution_unit_0_register_file_0_n_188));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_188),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_173 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[8]),.ZN(execution_unit_0_register_file_0_n_105_165));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_17 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_73_9));
	INV_X1_LVT execution_unit_0register_file_0i_73_18 (.A(execution_unit_0_register_file_0_n_73_9),.ZN(execution_unit_0_register_file_0_n_169));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_169),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_174 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[8]),.ZN(execution_unit_0_register_file_0_n_105_166));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_17 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_66_9));
	INV_X1_LVT execution_unit_0register_file_0i_66_18 (.A(execution_unit_0_register_file_0_n_66_9),.ZN(execution_unit_0_register_file_0_n_150));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_150),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_175 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[8]),.ZN(execution_unit_0_register_file_0_n_105_167));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_17 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_59_9));
	INV_X1_LVT execution_unit_0register_file_0i_59_18 (.A(execution_unit_0_register_file_0_n_59_9),.ZN(execution_unit_0_register_file_0_n_131));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_131),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_176 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[8]),.ZN(execution_unit_0_register_file_0_n_105_168));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_177 (.A1(execution_unit_0_register_file_0_n_105_165),.A2(execution_unit_0_register_file_0_n_105_166),.A3(execution_unit_0_register_file_0_n_105_167),.A4(execution_unit_0_register_file_0_n_105_168),.ZN(execution_unit_0_register_file_0_n_105_169));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_17 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_52_9));
	INV_X1_LVT execution_unit_0register_file_0i_52_18 (.A(execution_unit_0_register_file_0_n_52_9),.ZN(execution_unit_0_register_file_0_n_112));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_112),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_178 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[8]),.ZN(execution_unit_0_register_file_0_n_105_170));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_17 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_45_9));
	INV_X1_LVT execution_unit_0register_file_0i_45_18 (.A(execution_unit_0_register_file_0_n_45_9),.ZN(execution_unit_0_register_file_0_n_93));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_93),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_179 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[8]),.ZN(execution_unit_0_register_file_0_n_105_171));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_17 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_38_9));
	INV_X1_LVT execution_unit_0register_file_0i_38_18 (.A(execution_unit_0_register_file_0_n_38_9),.ZN(execution_unit_0_register_file_0_n_74));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_74),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_180 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[8]),.ZN(execution_unit_0_register_file_0_n_105_172));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_17 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_31_9));
	INV_X1_LVT execution_unit_0register_file_0i_31_18 (.A(execution_unit_0_register_file_0_n_31_9),.ZN(execution_unit_0_register_file_0_n_55));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_55),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_181 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[8]),.ZN(execution_unit_0_register_file_0_n_105_173));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_182 (.A1(execution_unit_0_register_file_0_n_105_170),.A2(execution_unit_0_register_file_0_n_105_171),.A3(execution_unit_0_register_file_0_n_105_172),.A4(execution_unit_0_register_file_0_n_105_173),.ZN(execution_unit_0_register_file_0_n_105_174));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_17 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_87_9));
	INV_X1_LVT execution_unit_0register_file_0i_87_18 (.A(execution_unit_0_register_file_0_n_87_9),.ZN(execution_unit_0_register_file_0_n_207));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_207),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[8]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_183 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[8]),.ZN(execution_unit_0_register_file_0_n_105_175));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_184 (.A1(execution_unit_0_register_file_0_n_105_164),.A2(execution_unit_0_register_file_0_n_105_169),.A3(execution_unit_0_register_file_0_n_105_174),.A4(execution_unit_0_register_file_0_n_105_175),.ZN(execution_unit_0_register_file_0_n_105_176));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_185 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[8]),.ZN(execution_unit_0_register_file_0_n_105_177));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_17 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_101_9));
	INV_X1_LVT execution_unit_0register_file_0i_101_18 (.A(execution_unit_0_register_file_0_n_101_9),.ZN(execution_unit_0_register_file_0_n_245));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_245),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_186 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[8]),.ZN(execution_unit_0_register_file_0_n_105_178));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_17 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[8]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(pc_sw[8]),.ZN(execution_unit_0_register_file_0_n_94_9));
	INV_X1_LVT execution_unit_0register_file_0i_94_18 (.A(execution_unit_0_register_file_0_n_94_9),.ZN(execution_unit_0_register_file_0_n_226));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b8___05F05d (.D(execution_unit_0_register_file_0_n_226),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[8]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_187 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[8]),.ZN(execution_unit_0_register_file_0_n_105_179));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_188 (.A1(execution_unit_0_register_file_0_n_105_176),.A2(execution_unit_0_register_file_0_n_105_177),.A3(execution_unit_0_register_file_0_n_105_178),.A4(execution_unit_0_register_file_0_n_105_179),.ZN(execution_unit_0_reg_src[8]));
	HA_X1_LVT execution_unit_0register_file_0i_106_7 (.A(execution_unit_0_reg_src[8]),.B(execution_unit_0_register_file_0_n_106_5),.CO(execution_unit_0_register_file_0_n_106_6),.S(execution_unit_0_register_file_0_n_262));
	HA_X1_LVT execution_unit_0register_file_0i_106_8 (.A(execution_unit_0_reg_src[9]),.B(execution_unit_0_register_file_0_n_106_6),.CO(execution_unit_0_register_file_0_n_106_7),.S(execution_unit_0_register_file_0_n_263));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_16 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(pc_sw[9]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[9]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_263),.ZN(execution_unit_0_register_file_0_n_109_8));
	INV_X1_LVT execution_unit_0register_file_0i_109_17 (.A(execution_unit_0_register_file_0_n_109_8),.ZN(execution_unit_0_register_file_0_n_281));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_281),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_192 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[9]),.ZN(execution_unit_0_register_file_0_n_105_183));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_193 (.A1(execution_unit_0_register_file_0_n_105_180),.A2(execution_unit_0_register_file_0_n_105_181),.A3(execution_unit_0_register_file_0_n_105_182),.A4(execution_unit_0_register_file_0_n_105_183),.ZN(execution_unit_0_register_file_0_n_105_184));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_19 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_80_10));
	INV_X1_LVT execution_unit_0register_file_0i_80_20 (.A(execution_unit_0_register_file_0_n_80_10),.ZN(execution_unit_0_register_file_0_n_189));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_189),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_194 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[9]),.ZN(execution_unit_0_register_file_0_n_105_185));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_19 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_73_10));
	INV_X1_LVT execution_unit_0register_file_0i_73_20 (.A(execution_unit_0_register_file_0_n_73_10),.ZN(execution_unit_0_register_file_0_n_170));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_170),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_195 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[9]),.ZN(execution_unit_0_register_file_0_n_105_186));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_19 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_66_10));
	INV_X1_LVT execution_unit_0register_file_0i_66_20 (.A(execution_unit_0_register_file_0_n_66_10),.ZN(execution_unit_0_register_file_0_n_151));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_151),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_196 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[9]),.ZN(execution_unit_0_register_file_0_n_105_187));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_19 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_59_10));
	INV_X1_LVT execution_unit_0register_file_0i_59_20 (.A(execution_unit_0_register_file_0_n_59_10),.ZN(execution_unit_0_register_file_0_n_132));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_132),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_197 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[9]),.ZN(execution_unit_0_register_file_0_n_105_188));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_198 (.A1(execution_unit_0_register_file_0_n_105_185),.A2(execution_unit_0_register_file_0_n_105_186),.A3(execution_unit_0_register_file_0_n_105_187),.A4(execution_unit_0_register_file_0_n_105_188),.ZN(execution_unit_0_register_file_0_n_105_189));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_19 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_52_10));
	INV_X1_LVT execution_unit_0register_file_0i_52_20 (.A(execution_unit_0_register_file_0_n_52_10),.ZN(execution_unit_0_register_file_0_n_113));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_113),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_199 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[9]),.ZN(execution_unit_0_register_file_0_n_105_190));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_19 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_45_10));
	INV_X1_LVT execution_unit_0register_file_0i_45_20 (.A(execution_unit_0_register_file_0_n_45_10),.ZN(execution_unit_0_register_file_0_n_94));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_94),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_200 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[9]),.ZN(execution_unit_0_register_file_0_n_105_191));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_19 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_38_10));
	INV_X1_LVT execution_unit_0register_file_0i_38_20 (.A(execution_unit_0_register_file_0_n_38_10),.ZN(execution_unit_0_register_file_0_n_75));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_75),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_201 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[9]),.ZN(execution_unit_0_register_file_0_n_105_192));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_19 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_31_10));
	INV_X1_LVT execution_unit_0register_file_0i_31_20 (.A(execution_unit_0_register_file_0_n_31_10),.ZN(execution_unit_0_register_file_0_n_56));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_56),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_202 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[9]),.ZN(execution_unit_0_register_file_0_n_105_193));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_203 (.A1(execution_unit_0_register_file_0_n_105_190),.A2(execution_unit_0_register_file_0_n_105_191),.A3(execution_unit_0_register_file_0_n_105_192),.A4(execution_unit_0_register_file_0_n_105_193),.ZN(execution_unit_0_register_file_0_n_105_194));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_19 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_87_10));
	INV_X1_LVT execution_unit_0register_file_0i_87_20 (.A(execution_unit_0_register_file_0_n_87_10),.ZN(execution_unit_0_register_file_0_n_208));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_208),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[9]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_204 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[9]),.ZN(execution_unit_0_register_file_0_n_105_195));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_205 (.A1(execution_unit_0_register_file_0_n_105_184),.A2(execution_unit_0_register_file_0_n_105_189),.A3(execution_unit_0_register_file_0_n_105_194),.A4(execution_unit_0_register_file_0_n_105_195),.ZN(execution_unit_0_register_file_0_n_105_196));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_206 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[9]),.ZN(execution_unit_0_register_file_0_n_105_197));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_19 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_101_10));
	INV_X1_LVT execution_unit_0register_file_0i_101_20 (.A(execution_unit_0_register_file_0_n_101_10),.ZN(execution_unit_0_register_file_0_n_246));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_246),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_207 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[9]),.ZN(execution_unit_0_register_file_0_n_105_198));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_19 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[9]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(pc_sw[9]),.ZN(execution_unit_0_register_file_0_n_94_10));
	INV_X1_LVT execution_unit_0register_file_0i_94_20 (.A(execution_unit_0_register_file_0_n_94_10),.ZN(execution_unit_0_register_file_0_n_227));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b9___05F05d (.D(execution_unit_0_register_file_0_n_227),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[9]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_208 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[9]),.ZN(execution_unit_0_register_file_0_n_105_199));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_209 (.A1(execution_unit_0_register_file_0_n_105_196),.A2(execution_unit_0_register_file_0_n_105_197),.A3(execution_unit_0_register_file_0_n_105_198),.A4(execution_unit_0_register_file_0_n_105_199),.ZN(execution_unit_0_reg_src[9]));
	HA_X1_LVT execution_unit_0register_file_0i_22_9 (.A(execution_unit_0_reg_src[9]),.B(execution_unit_0_register_file_0_n_22_8),.CO(execution_unit_0_register_file_0_n_22_9),.S(execution_unit_0_register_file_0_reg_incr_val[9]));
	HA_X1_LVT execution_unit_0register_file_0i_22_10 (.A(execution_unit_0_reg_src[10]),.B(execution_unit_0_register_file_0_n_22_9),.CO(execution_unit_0_register_file_0_n_22_10),.S(execution_unit_0_register_file_0_reg_incr_val[10]));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_21 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_24_11));
	INV_X1_LVT execution_unit_0register_file_0i_24_22 (.A(execution_unit_0_register_file_0_n_24_11),.ZN(execution_unit_0_register_file_0_n_38));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_38),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_210 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[10]),.ZN(execution_unit_0_register_file_0_n_105_200));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b10___05F05d (.D(pc_sw[10]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_211 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[10]),.ZN(execution_unit_0_register_file_0_n_105_201));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b10___05F05d (.D(1'b0),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_register_file_0_n_5),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_212 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_register_file_0_n_5),.ZN(execution_unit_0_register_file_0_n_105_202));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_18 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(pc_sw[10]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[10]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_264),.ZN(execution_unit_0_register_file_0_n_109_9));
	INV_X1_LVT execution_unit_0register_file_0i_109_19 (.A(execution_unit_0_register_file_0_n_109_9),.ZN(execution_unit_0_register_file_0_n_282));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_282),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_213 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[10]),.ZN(execution_unit_0_register_file_0_n_105_203));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_214 (.A1(execution_unit_0_register_file_0_n_105_200),.A2(execution_unit_0_register_file_0_n_105_201),.A3(execution_unit_0_register_file_0_n_105_202),.A4(execution_unit_0_register_file_0_n_105_203),.ZN(execution_unit_0_register_file_0_n_105_204));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_21 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_80_11));
	INV_X1_LVT execution_unit_0register_file_0i_80_22 (.A(execution_unit_0_register_file_0_n_80_11),.ZN(execution_unit_0_register_file_0_n_190));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_190),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_215 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[10]),.ZN(execution_unit_0_register_file_0_n_105_205));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_21 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_73_11));
	INV_X1_LVT execution_unit_0register_file_0i_73_22 (.A(execution_unit_0_register_file_0_n_73_11),.ZN(execution_unit_0_register_file_0_n_171));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_171),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_216 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[10]),.ZN(execution_unit_0_register_file_0_n_105_206));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_21 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_66_11));
	INV_X1_LVT execution_unit_0register_file_0i_66_22 (.A(execution_unit_0_register_file_0_n_66_11),.ZN(execution_unit_0_register_file_0_n_152));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_152),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_217 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[10]),.ZN(execution_unit_0_register_file_0_n_105_207));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_21 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_59_11));
	INV_X1_LVT execution_unit_0register_file_0i_59_22 (.A(execution_unit_0_register_file_0_n_59_11),.ZN(execution_unit_0_register_file_0_n_133));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_133),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_218 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[10]),.ZN(execution_unit_0_register_file_0_n_105_208));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_219 (.A1(execution_unit_0_register_file_0_n_105_205),.A2(execution_unit_0_register_file_0_n_105_206),.A3(execution_unit_0_register_file_0_n_105_207),.A4(execution_unit_0_register_file_0_n_105_208),.ZN(execution_unit_0_register_file_0_n_105_209));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_21 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_52_11));
	INV_X1_LVT execution_unit_0register_file_0i_52_22 (.A(execution_unit_0_register_file_0_n_52_11),.ZN(execution_unit_0_register_file_0_n_114));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_114),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_220 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[10]),.ZN(execution_unit_0_register_file_0_n_105_210));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_21 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_45_11));
	INV_X1_LVT execution_unit_0register_file_0i_45_22 (.A(execution_unit_0_register_file_0_n_45_11),.ZN(execution_unit_0_register_file_0_n_95));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_95),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_221 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[10]),.ZN(execution_unit_0_register_file_0_n_105_211));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_21 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_38_11));
	INV_X1_LVT execution_unit_0register_file_0i_38_22 (.A(execution_unit_0_register_file_0_n_38_11),.ZN(execution_unit_0_register_file_0_n_76));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_76),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_222 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[10]),.ZN(execution_unit_0_register_file_0_n_105_212));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_21 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_31_11));
	INV_X1_LVT execution_unit_0register_file_0i_31_22 (.A(execution_unit_0_register_file_0_n_31_11),.ZN(execution_unit_0_register_file_0_n_57));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_57),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_223 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[10]),.ZN(execution_unit_0_register_file_0_n_105_213));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_224 (.A1(execution_unit_0_register_file_0_n_105_210),.A2(execution_unit_0_register_file_0_n_105_211),.A3(execution_unit_0_register_file_0_n_105_212),.A4(execution_unit_0_register_file_0_n_105_213),.ZN(execution_unit_0_register_file_0_n_105_214));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_21 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_87_11));
	INV_X1_LVT execution_unit_0register_file_0i_87_22 (.A(execution_unit_0_register_file_0_n_87_11),.ZN(execution_unit_0_register_file_0_n_209));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_209),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[10]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_225 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[10]),.ZN(execution_unit_0_register_file_0_n_105_215));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_226 (.A1(execution_unit_0_register_file_0_n_105_204),.A2(execution_unit_0_register_file_0_n_105_209),.A3(execution_unit_0_register_file_0_n_105_214),.A4(execution_unit_0_register_file_0_n_105_215),.ZN(execution_unit_0_register_file_0_n_105_216));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_227 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[10]),.ZN(execution_unit_0_register_file_0_n_105_217));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_21 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_101_11));
	INV_X1_LVT execution_unit_0register_file_0i_101_22 (.A(execution_unit_0_register_file_0_n_101_11),.ZN(execution_unit_0_register_file_0_n_247));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_247),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_228 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[10]),.ZN(execution_unit_0_register_file_0_n_105_218));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_21 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[10]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(pc_sw[10]),.ZN(execution_unit_0_register_file_0_n_94_11));
	INV_X1_LVT execution_unit_0register_file_0i_94_22 (.A(execution_unit_0_register_file_0_n_94_11),.ZN(execution_unit_0_register_file_0_n_228));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b10___05F05d (.D(execution_unit_0_register_file_0_n_228),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[10]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_229 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[10]),.ZN(execution_unit_0_register_file_0_n_105_219));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_230 (.A1(execution_unit_0_register_file_0_n_105_216),.A2(execution_unit_0_register_file_0_n_105_217),.A3(execution_unit_0_register_file_0_n_105_218),.A4(execution_unit_0_register_file_0_n_105_219),.ZN(execution_unit_0_reg_src[10]));
	HA_X1_LVT execution_unit_0register_file_0i_106_9 (.A(execution_unit_0_reg_src[10]),.B(execution_unit_0_register_file_0_n_106_7),.CO(execution_unit_0_register_file_0_n_106_8),.S(execution_unit_0_register_file_0_n_264));
	HA_X1_LVT execution_unit_0register_file_0i_106_10 (.A(execution_unit_0_reg_src[11]),.B(execution_unit_0_register_file_0_n_106_8),.CO(execution_unit_0_register_file_0_n_106_9),.S(execution_unit_0_register_file_0_n_265));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_20 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(pc_sw[11]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[11]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_265),.ZN(execution_unit_0_register_file_0_n_109_10));
	INV_X1_LVT execution_unit_0register_file_0i_109_21 (.A(execution_unit_0_register_file_0_n_109_10),.ZN(execution_unit_0_register_file_0_n_283));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_283),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_234 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[11]),.ZN(execution_unit_0_register_file_0_n_105_223));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_235 (.A1(execution_unit_0_register_file_0_n_105_220),.A2(execution_unit_0_register_file_0_n_105_221),.A3(execution_unit_0_register_file_0_n_105_222),.A4(execution_unit_0_register_file_0_n_105_223),.ZN(execution_unit_0_register_file_0_n_105_224));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_23 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_80_12));
	INV_X1_LVT execution_unit_0register_file_0i_80_24 (.A(execution_unit_0_register_file_0_n_80_12),.ZN(execution_unit_0_register_file_0_n_191));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_191),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_236 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[11]),.ZN(execution_unit_0_register_file_0_n_105_225));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_23 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_73_12));
	INV_X1_LVT execution_unit_0register_file_0i_73_24 (.A(execution_unit_0_register_file_0_n_73_12),.ZN(execution_unit_0_register_file_0_n_172));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_172),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_237 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[11]),.ZN(execution_unit_0_register_file_0_n_105_226));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_23 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_66_12));
	INV_X1_LVT execution_unit_0register_file_0i_66_24 (.A(execution_unit_0_register_file_0_n_66_12),.ZN(execution_unit_0_register_file_0_n_153));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_153),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_238 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[11]),.ZN(execution_unit_0_register_file_0_n_105_227));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_23 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_59_12));
	INV_X1_LVT execution_unit_0register_file_0i_59_24 (.A(execution_unit_0_register_file_0_n_59_12),.ZN(execution_unit_0_register_file_0_n_134));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_134),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_239 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[11]),.ZN(execution_unit_0_register_file_0_n_105_228));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_240 (.A1(execution_unit_0_register_file_0_n_105_225),.A2(execution_unit_0_register_file_0_n_105_226),.A3(execution_unit_0_register_file_0_n_105_227),.A4(execution_unit_0_register_file_0_n_105_228),.ZN(execution_unit_0_register_file_0_n_105_229));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_23 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_52_12));
	INV_X1_LVT execution_unit_0register_file_0i_52_24 (.A(execution_unit_0_register_file_0_n_52_12),.ZN(execution_unit_0_register_file_0_n_115));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_115),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_241 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[11]),.ZN(execution_unit_0_register_file_0_n_105_230));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_23 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_45_12));
	INV_X1_LVT execution_unit_0register_file_0i_45_24 (.A(execution_unit_0_register_file_0_n_45_12),.ZN(execution_unit_0_register_file_0_n_96));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_96),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_242 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[11]),.ZN(execution_unit_0_register_file_0_n_105_231));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_23 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_38_12));
	INV_X1_LVT execution_unit_0register_file_0i_38_24 (.A(execution_unit_0_register_file_0_n_38_12),.ZN(execution_unit_0_register_file_0_n_77));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_77),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_243 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[11]),.ZN(execution_unit_0_register_file_0_n_105_232));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_23 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_31_12));
	INV_X1_LVT execution_unit_0register_file_0i_31_24 (.A(execution_unit_0_register_file_0_n_31_12),.ZN(execution_unit_0_register_file_0_n_58));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_58),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_244 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[11]),.ZN(execution_unit_0_register_file_0_n_105_233));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_245 (.A1(execution_unit_0_register_file_0_n_105_230),.A2(execution_unit_0_register_file_0_n_105_231),.A3(execution_unit_0_register_file_0_n_105_232),.A4(execution_unit_0_register_file_0_n_105_233),.ZN(execution_unit_0_register_file_0_n_105_234));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_23 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_87_12));
	INV_X1_LVT execution_unit_0register_file_0i_87_24 (.A(execution_unit_0_register_file_0_n_87_12),.ZN(execution_unit_0_register_file_0_n_210));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_210),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[11]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_246 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[11]),.ZN(execution_unit_0_register_file_0_n_105_235));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_247 (.A1(execution_unit_0_register_file_0_n_105_224),.A2(execution_unit_0_register_file_0_n_105_229),.A3(execution_unit_0_register_file_0_n_105_234),.A4(execution_unit_0_register_file_0_n_105_235),.ZN(execution_unit_0_register_file_0_n_105_236));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_248 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[11]),.ZN(execution_unit_0_register_file_0_n_105_237));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_23 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_101_12));
	INV_X1_LVT execution_unit_0register_file_0i_101_24 (.A(execution_unit_0_register_file_0_n_101_12),.ZN(execution_unit_0_register_file_0_n_248));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_248),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_249 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[11]),.ZN(execution_unit_0_register_file_0_n_105_238));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_23 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[11]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(pc_sw[11]),.ZN(execution_unit_0_register_file_0_n_94_12));
	INV_X1_LVT execution_unit_0register_file_0i_94_24 (.A(execution_unit_0_register_file_0_n_94_12),.ZN(execution_unit_0_register_file_0_n_229));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b11___05F05d (.D(execution_unit_0_register_file_0_n_229),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[11]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_250 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[11]),.ZN(execution_unit_0_register_file_0_n_105_239));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_251 (.A1(execution_unit_0_register_file_0_n_105_236),.A2(execution_unit_0_register_file_0_n_105_237),.A3(execution_unit_0_register_file_0_n_105_238),.A4(execution_unit_0_register_file_0_n_105_239),.ZN(execution_unit_0_reg_src[11]));
	HA_X1_LVT execution_unit_0register_file_0i_22_11 (.A(execution_unit_0_reg_src[11]),.B(execution_unit_0_register_file_0_n_22_10),.CO(execution_unit_0_register_file_0_n_22_11),.S(execution_unit_0_register_file_0_reg_incr_val[11]));
	HA_X1_LVT execution_unit_0register_file_0i_22_12 (.A(execution_unit_0_reg_src[12]),.B(execution_unit_0_register_file_0_n_22_11),.CO(execution_unit_0_register_file_0_n_22_12),.S(execution_unit_0_register_file_0_reg_incr_val[12]));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_25 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_24_13));
	INV_X1_LVT execution_unit_0register_file_0i_24_26 (.A(execution_unit_0_register_file_0_n_24_13),.ZN(execution_unit_0_register_file_0_n_40));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_40),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_252 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[12]),.ZN(execution_unit_0_register_file_0_n_105_240));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b12___05F05d (.D(pc_sw[12]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_253 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[12]),.ZN(execution_unit_0_register_file_0_n_105_241));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b12___05F05d (.D(1'b0),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_register_file_0_n_3),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_254 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_register_file_0_n_3),.ZN(execution_unit_0_register_file_0_n_105_242));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_22 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(pc_sw[12]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[12]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_266),.ZN(execution_unit_0_register_file_0_n_109_11));
	INV_X1_LVT execution_unit_0register_file_0i_109_23 (.A(execution_unit_0_register_file_0_n_109_11),.ZN(execution_unit_0_register_file_0_n_284));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_284),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_255 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[12]),.ZN(execution_unit_0_register_file_0_n_105_243));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_256 (.A1(execution_unit_0_register_file_0_n_105_240),.A2(execution_unit_0_register_file_0_n_105_241),.A3(execution_unit_0_register_file_0_n_105_242),.A4(execution_unit_0_register_file_0_n_105_243),.ZN(execution_unit_0_register_file_0_n_105_244));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_25 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_80_13));
	INV_X1_LVT execution_unit_0register_file_0i_80_26 (.A(execution_unit_0_register_file_0_n_80_13),.ZN(execution_unit_0_register_file_0_n_192));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_192),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_257 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[12]),.ZN(execution_unit_0_register_file_0_n_105_245));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_25 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_73_13));
	INV_X1_LVT execution_unit_0register_file_0i_73_26 (.A(execution_unit_0_register_file_0_n_73_13),.ZN(execution_unit_0_register_file_0_n_173));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_173),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_258 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[12]),.ZN(execution_unit_0_register_file_0_n_105_246));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_25 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_66_13));
	INV_X1_LVT execution_unit_0register_file_0i_66_26 (.A(execution_unit_0_register_file_0_n_66_13),.ZN(execution_unit_0_register_file_0_n_154));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_154),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_259 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[12]),.ZN(execution_unit_0_register_file_0_n_105_247));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_25 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_59_13));
	INV_X1_LVT execution_unit_0register_file_0i_59_26 (.A(execution_unit_0_register_file_0_n_59_13),.ZN(execution_unit_0_register_file_0_n_135));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_135),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_260 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[12]),.ZN(execution_unit_0_register_file_0_n_105_248));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_261 (.A1(execution_unit_0_register_file_0_n_105_245),.A2(execution_unit_0_register_file_0_n_105_246),.A3(execution_unit_0_register_file_0_n_105_247),.A4(execution_unit_0_register_file_0_n_105_248),.ZN(execution_unit_0_register_file_0_n_105_249));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_25 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_52_13));
	INV_X1_LVT execution_unit_0register_file_0i_52_26 (.A(execution_unit_0_register_file_0_n_52_13),.ZN(execution_unit_0_register_file_0_n_116));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_116),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_262 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[12]),.ZN(execution_unit_0_register_file_0_n_105_250));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_25 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_45_13));
	INV_X1_LVT execution_unit_0register_file_0i_45_26 (.A(execution_unit_0_register_file_0_n_45_13),.ZN(execution_unit_0_register_file_0_n_97));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_97),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_263 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[12]),.ZN(execution_unit_0_register_file_0_n_105_251));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_25 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_38_13));
	INV_X1_LVT execution_unit_0register_file_0i_38_26 (.A(execution_unit_0_register_file_0_n_38_13),.ZN(execution_unit_0_register_file_0_n_78));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_78),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_264 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[12]),.ZN(execution_unit_0_register_file_0_n_105_252));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_25 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_31_13));
	INV_X1_LVT execution_unit_0register_file_0i_31_26 (.A(execution_unit_0_register_file_0_n_31_13),.ZN(execution_unit_0_register_file_0_n_59));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_59),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_265 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[12]),.ZN(execution_unit_0_register_file_0_n_105_253));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_266 (.A1(execution_unit_0_register_file_0_n_105_250),.A2(execution_unit_0_register_file_0_n_105_251),.A3(execution_unit_0_register_file_0_n_105_252),.A4(execution_unit_0_register_file_0_n_105_253),.ZN(execution_unit_0_register_file_0_n_105_254));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_25 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_87_13));
	INV_X1_LVT execution_unit_0register_file_0i_87_26 (.A(execution_unit_0_register_file_0_n_87_13),.ZN(execution_unit_0_register_file_0_n_211));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_211),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[12]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_267 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[12]),.ZN(execution_unit_0_register_file_0_n_105_255));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_268 (.A1(execution_unit_0_register_file_0_n_105_244),.A2(execution_unit_0_register_file_0_n_105_249),.A3(execution_unit_0_register_file_0_n_105_254),.A4(execution_unit_0_register_file_0_n_105_255),.ZN(execution_unit_0_register_file_0_n_105_256));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_269 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[12]),.ZN(execution_unit_0_register_file_0_n_105_257));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_25 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_101_13));
	INV_X1_LVT execution_unit_0register_file_0i_101_26 (.A(execution_unit_0_register_file_0_n_101_13),.ZN(execution_unit_0_register_file_0_n_249));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_249),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_270 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[12]),.ZN(execution_unit_0_register_file_0_n_105_258));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_25 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[12]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(pc_sw[12]),.ZN(execution_unit_0_register_file_0_n_94_13));
	INV_X1_LVT execution_unit_0register_file_0i_94_26 (.A(execution_unit_0_register_file_0_n_94_13),.ZN(execution_unit_0_register_file_0_n_230));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b12___05F05d (.D(execution_unit_0_register_file_0_n_230),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[12]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_271 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[12]),.ZN(execution_unit_0_register_file_0_n_105_259));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_272 (.A1(execution_unit_0_register_file_0_n_105_256),.A2(execution_unit_0_register_file_0_n_105_257),.A3(execution_unit_0_register_file_0_n_105_258),.A4(execution_unit_0_register_file_0_n_105_259),.ZN(execution_unit_0_reg_src[12]));
	HA_X1_LVT execution_unit_0register_file_0i_106_11 (.A(execution_unit_0_reg_src[12]),.B(execution_unit_0_register_file_0_n_106_9),.CO(execution_unit_0_register_file_0_n_106_10),.S(execution_unit_0_register_file_0_n_266));
	HA_X1_LVT execution_unit_0register_file_0i_106_12 (.A(execution_unit_0_reg_src[13]),.B(execution_unit_0_register_file_0_n_106_10),.CO(execution_unit_0_register_file_0_n_106_11),.S(execution_unit_0_register_file_0_n_267));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_24 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(pc_sw[13]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[13]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_267),.ZN(execution_unit_0_register_file_0_n_109_12));
	INV_X1_LVT execution_unit_0register_file_0i_109_25 (.A(execution_unit_0_register_file_0_n_109_12),.ZN(execution_unit_0_register_file_0_n_285));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_285),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_276 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[13]),.ZN(execution_unit_0_register_file_0_n_105_263));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_277 (.A1(execution_unit_0_register_file_0_n_105_260),.A2(execution_unit_0_register_file_0_n_105_261),.A3(execution_unit_0_register_file_0_n_105_262),.A4(execution_unit_0_register_file_0_n_105_263),.ZN(execution_unit_0_register_file_0_n_105_264));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_27 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_80_14));
	INV_X1_LVT execution_unit_0register_file_0i_80_28 (.A(execution_unit_0_register_file_0_n_80_14),.ZN(execution_unit_0_register_file_0_n_193));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_193),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_278 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[13]),.ZN(execution_unit_0_register_file_0_n_105_265));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_27 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_73_14));
	INV_X1_LVT execution_unit_0register_file_0i_73_28 (.A(execution_unit_0_register_file_0_n_73_14),.ZN(execution_unit_0_register_file_0_n_174));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_174),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_279 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[13]),.ZN(execution_unit_0_register_file_0_n_105_266));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_27 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_66_14));
	INV_X1_LVT execution_unit_0register_file_0i_66_28 (.A(execution_unit_0_register_file_0_n_66_14),.ZN(execution_unit_0_register_file_0_n_155));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_155),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_280 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[13]),.ZN(execution_unit_0_register_file_0_n_105_267));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_27 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_59_14));
	INV_X1_LVT execution_unit_0register_file_0i_59_28 (.A(execution_unit_0_register_file_0_n_59_14),.ZN(execution_unit_0_register_file_0_n_136));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_136),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_281 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[13]),.ZN(execution_unit_0_register_file_0_n_105_268));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_282 (.A1(execution_unit_0_register_file_0_n_105_265),.A2(execution_unit_0_register_file_0_n_105_266),.A3(execution_unit_0_register_file_0_n_105_267),.A4(execution_unit_0_register_file_0_n_105_268),.ZN(execution_unit_0_register_file_0_n_105_269));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_27 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_52_14));
	INV_X1_LVT execution_unit_0register_file_0i_52_28 (.A(execution_unit_0_register_file_0_n_52_14),.ZN(execution_unit_0_register_file_0_n_117));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_117),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_283 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[13]),.ZN(execution_unit_0_register_file_0_n_105_270));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_27 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_45_14));
	INV_X1_LVT execution_unit_0register_file_0i_45_28 (.A(execution_unit_0_register_file_0_n_45_14),.ZN(execution_unit_0_register_file_0_n_98));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_98),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_284 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[13]),.ZN(execution_unit_0_register_file_0_n_105_271));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_27 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_38_14));
	INV_X1_LVT execution_unit_0register_file_0i_38_28 (.A(execution_unit_0_register_file_0_n_38_14),.ZN(execution_unit_0_register_file_0_n_79));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_79),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_285 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[13]),.ZN(execution_unit_0_register_file_0_n_105_272));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_27 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_31_14));
	INV_X1_LVT execution_unit_0register_file_0i_31_28 (.A(execution_unit_0_register_file_0_n_31_14),.ZN(execution_unit_0_register_file_0_n_60));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_60),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_286 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[13]),.ZN(execution_unit_0_register_file_0_n_105_273));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_287 (.A1(execution_unit_0_register_file_0_n_105_270),.A2(execution_unit_0_register_file_0_n_105_271),.A3(execution_unit_0_register_file_0_n_105_272),.A4(execution_unit_0_register_file_0_n_105_273),.ZN(execution_unit_0_register_file_0_n_105_274));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_27 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_87_14));
	INV_X1_LVT execution_unit_0register_file_0i_87_28 (.A(execution_unit_0_register_file_0_n_87_14),.ZN(execution_unit_0_register_file_0_n_212));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_212),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[13]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_288 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[13]),.ZN(execution_unit_0_register_file_0_n_105_275));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_289 (.A1(execution_unit_0_register_file_0_n_105_264),.A2(execution_unit_0_register_file_0_n_105_269),.A3(execution_unit_0_register_file_0_n_105_274),.A4(execution_unit_0_register_file_0_n_105_275),.ZN(execution_unit_0_register_file_0_n_105_276));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_290 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[13]),.ZN(execution_unit_0_register_file_0_n_105_277));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_27 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_101_14));
	INV_X1_LVT execution_unit_0register_file_0i_101_28 (.A(execution_unit_0_register_file_0_n_101_14),.ZN(execution_unit_0_register_file_0_n_250));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_250),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_291 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[13]),.ZN(execution_unit_0_register_file_0_n_105_278));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_27 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[13]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(pc_sw[13]),.ZN(execution_unit_0_register_file_0_n_94_14));
	INV_X1_LVT execution_unit_0register_file_0i_94_28 (.A(execution_unit_0_register_file_0_n_94_14),.ZN(execution_unit_0_register_file_0_n_231));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b13___05F05d (.D(execution_unit_0_register_file_0_n_231),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[13]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_292 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[13]),.ZN(execution_unit_0_register_file_0_n_105_279));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_293 (.A1(execution_unit_0_register_file_0_n_105_276),.A2(execution_unit_0_register_file_0_n_105_277),.A3(execution_unit_0_register_file_0_n_105_278),.A4(execution_unit_0_register_file_0_n_105_279),.ZN(execution_unit_0_reg_src[13]));
	HA_X1_LVT execution_unit_0register_file_0i_22_13 (.A(execution_unit_0_reg_src[13]),.B(execution_unit_0_register_file_0_n_22_12),.CO(execution_unit_0_register_file_0_n_22_13),.S(execution_unit_0_register_file_0_reg_incr_val[13]));
	HA_X1_LVT execution_unit_0register_file_0i_22_14 (.A(execution_unit_0_reg_src[14]),.B(execution_unit_0_register_file_0_n_22_13),.CO(execution_unit_0_register_file_0_n_22_14),.S(execution_unit_0_register_file_0_reg_incr_val[14]));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_29 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_24_15));
	INV_X1_LVT execution_unit_0register_file_0i_24_30 (.A(execution_unit_0_register_file_0_n_24_15),.ZN(execution_unit_0_register_file_0_n_42));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_42),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_294 (.A1(execution_unit_0_register_file_0_n_24),.A2(execution_unit_0_register_file_0_r4[14]),.ZN(execution_unit_0_register_file_0_n_105_280));
	DFFR_X1_LVT execution_unit_0register_file_0r3_reg___05F05b14___05F05d (.D(pc_sw[14]),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_23),.Q(execution_unit_0_register_file_0_r3[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_295 (.A1(execution_unit_0_register_file_0_n_22),.A2(execution_unit_0_register_file_0_r3[14]),.ZN(execution_unit_0_register_file_0_n_105_281));
	DFFR_X1_LVT execution_unit_0register_file_0r2_reg___05F05b14___05F05d (.D(1'b0),.RN(execution_unit_0_register_file_0_n_8),.CK(cpu_mclk),.Q(execution_unit_0_register_file_0_n_1),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_296 (.A1(execution_unit_0_register_file_0_n_21),.A2(execution_unit_0_register_file_0_n_1),.ZN(execution_unit_0_register_file_0_n_105_282));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_26 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(pc_sw[14]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[14]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_268),.ZN(execution_unit_0_register_file_0_n_109_13));
	INV_X1_LVT execution_unit_0register_file_0i_109_27 (.A(execution_unit_0_register_file_0_n_109_13),.ZN(execution_unit_0_register_file_0_n_286));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_286),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_297 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[14]),.ZN(execution_unit_0_register_file_0_n_105_283));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_298 (.A1(execution_unit_0_register_file_0_n_105_280),.A2(execution_unit_0_register_file_0_n_105_281),.A3(execution_unit_0_register_file_0_n_105_282),.A4(execution_unit_0_register_file_0_n_105_283),.ZN(execution_unit_0_register_file_0_n_105_284));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_29 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_80_15));
	INV_X1_LVT execution_unit_0register_file_0i_80_30 (.A(execution_unit_0_register_file_0_n_80_15),.ZN(execution_unit_0_register_file_0_n_194));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_194),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_299 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[14]),.ZN(execution_unit_0_register_file_0_n_105_285));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_29 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_73_15));
	INV_X1_LVT execution_unit_0register_file_0i_73_30 (.A(execution_unit_0_register_file_0_n_73_15),.ZN(execution_unit_0_register_file_0_n_175));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_175),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_300 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[14]),.ZN(execution_unit_0_register_file_0_n_105_286));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_29 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_66_15));
	INV_X1_LVT execution_unit_0register_file_0i_66_30 (.A(execution_unit_0_register_file_0_n_66_15),.ZN(execution_unit_0_register_file_0_n_156));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_156),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_301 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[14]),.ZN(execution_unit_0_register_file_0_n_105_287));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_29 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_59_15));
	INV_X1_LVT execution_unit_0register_file_0i_59_30 (.A(execution_unit_0_register_file_0_n_59_15),.ZN(execution_unit_0_register_file_0_n_137));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_137),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_302 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[14]),.ZN(execution_unit_0_register_file_0_n_105_288));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_303 (.A1(execution_unit_0_register_file_0_n_105_285),.A2(execution_unit_0_register_file_0_n_105_286),.A3(execution_unit_0_register_file_0_n_105_287),.A4(execution_unit_0_register_file_0_n_105_288),.ZN(execution_unit_0_register_file_0_n_105_289));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_29 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_52_15));
	INV_X1_LVT execution_unit_0register_file_0i_52_30 (.A(execution_unit_0_register_file_0_n_52_15),.ZN(execution_unit_0_register_file_0_n_118));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_118),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_304 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[14]),.ZN(execution_unit_0_register_file_0_n_105_290));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_29 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_45_15));
	INV_X1_LVT execution_unit_0register_file_0i_45_30 (.A(execution_unit_0_register_file_0_n_45_15),.ZN(execution_unit_0_register_file_0_n_99));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_99),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_305 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[14]),.ZN(execution_unit_0_register_file_0_n_105_291));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_29 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_38_15));
	INV_X1_LVT execution_unit_0register_file_0i_38_30 (.A(execution_unit_0_register_file_0_n_38_15),.ZN(execution_unit_0_register_file_0_n_80));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_80),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_306 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[14]),.ZN(execution_unit_0_register_file_0_n_105_292));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_29 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_31_15));
	INV_X1_LVT execution_unit_0register_file_0i_31_30 (.A(execution_unit_0_register_file_0_n_31_15),.ZN(execution_unit_0_register_file_0_n_61));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_61),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_307 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[14]),.ZN(execution_unit_0_register_file_0_n_105_293));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_308 (.A1(execution_unit_0_register_file_0_n_105_290),.A2(execution_unit_0_register_file_0_n_105_291),.A3(execution_unit_0_register_file_0_n_105_292),.A4(execution_unit_0_register_file_0_n_105_293),.ZN(execution_unit_0_register_file_0_n_105_294));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_29 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_87_15));
	INV_X1_LVT execution_unit_0register_file_0i_87_30 (.A(execution_unit_0_register_file_0_n_87_15),.ZN(execution_unit_0_register_file_0_n_213));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_213),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[14]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_309 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[14]),.ZN(execution_unit_0_register_file_0_n_105_295));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_310 (.A1(execution_unit_0_register_file_0_n_105_284),.A2(execution_unit_0_register_file_0_n_105_289),.A3(execution_unit_0_register_file_0_n_105_294),.A4(execution_unit_0_register_file_0_n_105_295),.ZN(execution_unit_0_register_file_0_n_105_296));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_311 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[14]),.ZN(execution_unit_0_register_file_0_n_105_297));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_29 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_101_15));
	INV_X1_LVT execution_unit_0register_file_0i_101_30 (.A(execution_unit_0_register_file_0_n_101_15),.ZN(execution_unit_0_register_file_0_n_251));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_251),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_312 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[14]),.ZN(execution_unit_0_register_file_0_n_105_298));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_29 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[14]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(pc_sw[14]),.ZN(execution_unit_0_register_file_0_n_94_15));
	INV_X1_LVT execution_unit_0register_file_0i_94_30 (.A(execution_unit_0_register_file_0_n_94_15),.ZN(execution_unit_0_register_file_0_n_232));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b14___05F05d (.D(execution_unit_0_register_file_0_n_232),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[14]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_313 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[14]),.ZN(execution_unit_0_register_file_0_n_105_299));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_314 (.A1(execution_unit_0_register_file_0_n_105_296),.A2(execution_unit_0_register_file_0_n_105_297),.A3(execution_unit_0_register_file_0_n_105_298),.A4(execution_unit_0_register_file_0_n_105_299),.ZN(execution_unit_0_reg_src[14]));
	HA_X1_LVT execution_unit_0register_file_0i_106_13 (.A(execution_unit_0_reg_src[14]),.B(execution_unit_0_register_file_0_n_106_11),.CO(execution_unit_0_register_file_0_n_106_12),.S(execution_unit_0_register_file_0_n_268));
	XNOR2_X1_LVT execution_unit_0register_file_0i_106_14 (.A(execution_unit_0_reg_src[15]),.B(execution_unit_0_register_file_0_n_106_12),.ZN(execution_unit_0_register_file_0_n_106_13));
	INV_X1_LVT execution_unit_0register_file_0i_106_15 (.A(execution_unit_0_register_file_0_n_106_13),.ZN(execution_unit_0_register_file_0_n_269));
	AOI222_X1_LVT execution_unit_0register_file_0i_109_28 (.A1(execution_unit_0_register_file_0_r1_wr),.A2(pc_sw[15]),.B1(execution_unit_0_register_file_0_n_272),.B2(eu_mab[15]),.C1(execution_unit_0_register_file_0_n_271),.C2(execution_unit_0_register_file_0_n_269),.ZN(execution_unit_0_register_file_0_n_109_14));
	INV_X1_LVT execution_unit_0register_file_0i_109_29 (.A(execution_unit_0_register_file_0_n_109_14),.ZN(execution_unit_0_register_file_0_n_287));
	DFFR_X1_LVT execution_unit_0register_file_0r1_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_287),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_270),.Q(execution_unit_0_register_file_0_r1[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_318 (.A1(execution_unit_0_register_file_0_inst_src_in),.A2(execution_unit_0_register_file_0_r1[15]),.ZN(execution_unit_0_register_file_0_n_105_303));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_319 (.A1(execution_unit_0_register_file_0_n_105_300),.A2(execution_unit_0_register_file_0_n_105_301),.A3(execution_unit_0_register_file_0_n_105_302),.A4(execution_unit_0_register_file_0_n_105_303),.ZN(execution_unit_0_register_file_0_n_105_304));
	AOI22_X1_LVT execution_unit_0register_file_0i_80_31 (.A1(execution_unit_0_register_file_0_n_80_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r12_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_80_16));
	INV_X1_LVT execution_unit_0register_file_0i_80_32 (.A(execution_unit_0_register_file_0_n_80_16),.ZN(execution_unit_0_register_file_0_n_195));
	DFFR_X1_LVT execution_unit_0register_file_0r12_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_195),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_179),.Q(execution_unit_0_register_file_0_r12[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_320 (.A1(execution_unit_0_register_file_0_n_178),.A2(execution_unit_0_register_file_0_r12[15]),.ZN(execution_unit_0_register_file_0_n_105_305));
	AOI22_X1_LVT execution_unit_0register_file_0i_73_31 (.A1(execution_unit_0_register_file_0_n_73_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r11_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_73_16));
	INV_X1_LVT execution_unit_0register_file_0i_73_32 (.A(execution_unit_0_register_file_0_n_73_16),.ZN(execution_unit_0_register_file_0_n_176));
	DFFR_X1_LVT execution_unit_0register_file_0r11_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_176),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_160),.Q(execution_unit_0_register_file_0_r11[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_321 (.A1(execution_unit_0_register_file_0_n_159),.A2(execution_unit_0_register_file_0_r11[15]),.ZN(execution_unit_0_register_file_0_n_105_306));
	AOI22_X1_LVT execution_unit_0register_file_0i_66_31 (.A1(execution_unit_0_register_file_0_n_66_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r10_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_66_16));
	INV_X1_LVT execution_unit_0register_file_0i_66_32 (.A(execution_unit_0_register_file_0_n_66_16),.ZN(execution_unit_0_register_file_0_n_157));
	DFFR_X1_LVT execution_unit_0register_file_0r10_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_157),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_141),.Q(execution_unit_0_register_file_0_r10[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_322 (.A1(execution_unit_0_register_file_0_n_140),.A2(execution_unit_0_register_file_0_r10[15]),.ZN(execution_unit_0_register_file_0_n_105_307));
	AOI22_X1_LVT execution_unit_0register_file_0i_59_31 (.A1(execution_unit_0_register_file_0_n_59_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r9_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_59_16));
	INV_X1_LVT execution_unit_0register_file_0i_59_32 (.A(execution_unit_0_register_file_0_n_59_16),.ZN(execution_unit_0_register_file_0_n_138));
	DFFR_X1_LVT execution_unit_0register_file_0r9_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_138),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_122),.Q(execution_unit_0_register_file_0_r9[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_323 (.A1(execution_unit_0_register_file_0_n_121),.A2(execution_unit_0_register_file_0_r9[15]),.ZN(execution_unit_0_register_file_0_n_105_308));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_324 (.A1(execution_unit_0_register_file_0_n_105_305),.A2(execution_unit_0_register_file_0_n_105_306),.A3(execution_unit_0_register_file_0_n_105_307),.A4(execution_unit_0_register_file_0_n_105_308),.ZN(execution_unit_0_register_file_0_n_105_309));
	AOI22_X1_LVT execution_unit_0register_file_0i_52_31 (.A1(execution_unit_0_register_file_0_n_52_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r8_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_52_16));
	INV_X1_LVT execution_unit_0register_file_0i_52_32 (.A(execution_unit_0_register_file_0_n_52_16),.ZN(execution_unit_0_register_file_0_n_119));
	DFFR_X1_LVT execution_unit_0register_file_0r8_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_119),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_103),.Q(execution_unit_0_register_file_0_r8[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_325 (.A1(execution_unit_0_register_file_0_n_102),.A2(execution_unit_0_register_file_0_r8[15]),.ZN(execution_unit_0_register_file_0_n_105_310));
	AOI22_X1_LVT execution_unit_0register_file_0i_45_31 (.A1(execution_unit_0_register_file_0_n_45_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r7_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_45_16));
	INV_X1_LVT execution_unit_0register_file_0i_45_32 (.A(execution_unit_0_register_file_0_n_45_16),.ZN(execution_unit_0_register_file_0_n_100));
	DFFR_X1_LVT execution_unit_0register_file_0r7_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_100),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_84),.Q(execution_unit_0_register_file_0_r7[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_326 (.A1(execution_unit_0_register_file_0_n_83),.A2(execution_unit_0_register_file_0_r7[15]),.ZN(execution_unit_0_register_file_0_n_105_311));
	AOI22_X1_LVT execution_unit_0register_file_0i_38_31 (.A1(execution_unit_0_register_file_0_n_38_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r6_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_38_16));
	INV_X1_LVT execution_unit_0register_file_0i_38_32 (.A(execution_unit_0_register_file_0_n_38_16),.ZN(execution_unit_0_register_file_0_n_81));
	DFFR_X1_LVT execution_unit_0register_file_0r6_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_81),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_65),.Q(execution_unit_0_register_file_0_r6[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_327 (.A1(execution_unit_0_register_file_0_n_64),.A2(execution_unit_0_register_file_0_r6[15]),.ZN(execution_unit_0_register_file_0_n_105_312));
	AOI22_X1_LVT execution_unit_0register_file_0i_31_31 (.A1(execution_unit_0_register_file_0_n_31_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r5_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_31_16));
	INV_X1_LVT execution_unit_0register_file_0i_31_32 (.A(execution_unit_0_register_file_0_n_31_16),.ZN(execution_unit_0_register_file_0_n_62));
	DFFR_X1_LVT execution_unit_0register_file_0r5_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_62),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_46),.Q(execution_unit_0_register_file_0_r5[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_328 (.A1(execution_unit_0_register_file_0_n_45),.A2(execution_unit_0_register_file_0_r5[15]),.ZN(execution_unit_0_register_file_0_n_105_313));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_329 (.A1(execution_unit_0_register_file_0_n_105_310),.A2(execution_unit_0_register_file_0_n_105_311),.A3(execution_unit_0_register_file_0_n_105_312),.A4(execution_unit_0_register_file_0_n_105_313),.ZN(execution_unit_0_register_file_0_n_105_314));
	AOI22_X1_LVT execution_unit_0register_file_0i_87_31 (.A1(execution_unit_0_register_file_0_n_87_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r13_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_87_16));
	INV_X1_LVT execution_unit_0register_file_0i_87_32 (.A(execution_unit_0_register_file_0_n_87_16),.ZN(execution_unit_0_register_file_0_n_214));
	DFFR_X1_LVT execution_unit_0register_file_0r13_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_214),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_198),.Q(execution_unit_0_register_file_0_r13[15]),.QN());
	AND2_X1_LVT execution_unit_0register_file_0i_105_330 (.A1(execution_unit_0_register_file_0_n_197),.A2(execution_unit_0_register_file_0_r13[15]),.ZN(execution_unit_0_register_file_0_n_105_315));
	NOR4_X1_LVT execution_unit_0register_file_0i_105_331 (.A1(execution_unit_0_register_file_0_n_105_304),.A2(execution_unit_0_register_file_0_n_105_309),.A3(execution_unit_0_register_file_0_n_105_314),.A4(execution_unit_0_register_file_0_n_105_315),.ZN(execution_unit_0_register_file_0_n_105_316));
	NAND2_X1_LVT execution_unit_0register_file_0i_105_332 (.A1(execution_unit_0_register_file_0_n_254),.A2(pc[15]),.ZN(execution_unit_0_register_file_0_n_105_317));
	AOI22_X1_LVT execution_unit_0register_file_0i_101_31 (.A1(execution_unit_0_register_file_0_n_101_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r15_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_101_16));
	INV_X1_LVT execution_unit_0register_file_0i_101_32 (.A(execution_unit_0_register_file_0_n_101_16),.ZN(execution_unit_0_register_file_0_n_252));
	DFFR_X1_LVT execution_unit_0register_file_0r15_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_252),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_236),.Q(execution_unit_0_register_file_0_r15[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_333 (.A1(execution_unit_0_register_file_0_n_235),.A2(execution_unit_0_register_file_0_r15[15]),.ZN(execution_unit_0_register_file_0_n_105_318));
	AOI22_X1_LVT execution_unit_0register_file_0i_94_31 (.A1(execution_unit_0_register_file_0_n_94_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r14_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_94_16));
	INV_X1_LVT execution_unit_0register_file_0i_94_32 (.A(execution_unit_0_register_file_0_n_94_16),.ZN(execution_unit_0_register_file_0_n_233));
	DFFR_X1_LVT execution_unit_0register_file_0r14_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_233),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_217),.Q(execution_unit_0_register_file_0_r14[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_105_334 (.A1(execution_unit_0_register_file_0_n_216),.A2(execution_unit_0_register_file_0_r14[15]),.ZN(execution_unit_0_register_file_0_n_105_319));
	NAND4_X1_LVT execution_unit_0register_file_0i_105_335 (.A1(execution_unit_0_register_file_0_n_105_316),.A2(execution_unit_0_register_file_0_n_105_317),.A3(execution_unit_0_register_file_0_n_105_318),.A4(execution_unit_0_register_file_0_n_105_319),.ZN(execution_unit_0_reg_src[15]));
	XNOR2_X1_LVT execution_unit_0register_file_0i_22_15 (.A(execution_unit_0_reg_src[15]),.B(execution_unit_0_register_file_0_n_22_14),.ZN(execution_unit_0_register_file_0_n_22_15));
	INV_X1_LVT execution_unit_0register_file_0i_22_16 (.A(execution_unit_0_register_file_0_n_22_15),.ZN(execution_unit_0_register_file_0_reg_incr_val[15]));
	AOI22_X1_LVT execution_unit_0register_file_0i_24_31 (.A1(execution_unit_0_register_file_0_n_24_0),.A2(execution_unit_0_register_file_0_reg_incr_val[15]),.B1(execution_unit_0_register_file_0_r4_wr),.B2(pc_sw[15]),.ZN(execution_unit_0_register_file_0_n_24_16));
	INV_X1_LVT execution_unit_0register_file_0i_24_32 (.A(execution_unit_0_register_file_0_n_24_16),.ZN(execution_unit_0_register_file_0_n_43));
	DFFR_X1_LVT execution_unit_0register_file_0r4_reg___05F05b15___05F05d (.D(execution_unit_0_register_file_0_n_43),.RN(execution_unit_0_register_file_0_n_8),.CK(execution_unit_0_register_file_0_n_27),.Q(execution_unit_0_register_file_0_r4[15]),.QN());
	NAND2_X1_LVT execution_unit_0register_file_0i_112_315 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[15]),.ZN(execution_unit_0_register_file_0_n_112_300));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_316 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[15]),.ZN(execution_unit_0_register_file_0_n_112_301));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_317 (.A1(inst_dest[2]),.A2(execution_unit_0_register_file_0_n_0),.ZN(execution_unit_0_register_file_0_n_112_302));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_318 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[15]),.ZN(execution_unit_0_register_file_0_n_112_303));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_319 (.A1(execution_unit_0_register_file_0_n_112_300),.A2(execution_unit_0_register_file_0_n_112_301),.A3(execution_unit_0_register_file_0_n_112_302),.A4(execution_unit_0_register_file_0_n_112_303),.ZN(execution_unit_0_register_file_0_n_112_304));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_320 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[15]),.ZN(execution_unit_0_register_file_0_n_112_305));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_321 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[15]),.ZN(execution_unit_0_register_file_0_n_112_306));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_322 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[15]),.ZN(execution_unit_0_register_file_0_n_112_307));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_323 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[15]),.ZN(execution_unit_0_register_file_0_n_112_308));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_324 (.A1(execution_unit_0_register_file_0_n_112_305),.A2(execution_unit_0_register_file_0_n_112_306),.A3(execution_unit_0_register_file_0_n_112_307),.A4(execution_unit_0_register_file_0_n_112_308),.ZN(execution_unit_0_register_file_0_n_112_309));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_325 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[15]),.ZN(execution_unit_0_register_file_0_n_112_310));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_326 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[15]),.ZN(execution_unit_0_register_file_0_n_112_311));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_327 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[15]),.ZN(execution_unit_0_register_file_0_n_112_312));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_328 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[15]),.ZN(execution_unit_0_register_file_0_n_112_313));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_329 (.A1(execution_unit_0_register_file_0_n_112_310),.A2(execution_unit_0_register_file_0_n_112_311),.A3(execution_unit_0_register_file_0_n_112_312),.A4(execution_unit_0_register_file_0_n_112_313),.ZN(execution_unit_0_register_file_0_n_112_314));
	AND2_X1_LVT execution_unit_0register_file_0i_112_330 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[15]),.ZN(execution_unit_0_register_file_0_n_112_315));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_331 (.A1(execution_unit_0_register_file_0_n_112_304),.A2(execution_unit_0_register_file_0_n_112_309),.A3(execution_unit_0_register_file_0_n_112_314),.A4(execution_unit_0_register_file_0_n_112_315),.ZN(execution_unit_0_register_file_0_n_112_316));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_332 (.A1(inst_dest[0]),.A2(pc[15]),.ZN(execution_unit_0_register_file_0_n_112_317));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_333 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[15]),.ZN(execution_unit_0_register_file_0_n_112_318));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_334 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[15]),.ZN(execution_unit_0_register_file_0_n_112_319));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_335 (.A1(execution_unit_0_register_file_0_n_112_316),.A2(execution_unit_0_register_file_0_n_112_317),.A3(execution_unit_0_register_file_0_n_112_318),.A4(execution_unit_0_register_file_0_n_112_319),.ZN(dbg_reg_din[15]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_294 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[14]),.ZN(execution_unit_0_register_file_0_n_112_280));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_295 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[14]),.ZN(execution_unit_0_register_file_0_n_112_281));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_296 (.A1(inst_dest[2]),.A2(execution_unit_0_register_file_0_n_1),.ZN(execution_unit_0_register_file_0_n_112_282));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_297 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[14]),.ZN(execution_unit_0_register_file_0_n_112_283));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_298 (.A1(execution_unit_0_register_file_0_n_112_280),.A2(execution_unit_0_register_file_0_n_112_281),.A3(execution_unit_0_register_file_0_n_112_282),.A4(execution_unit_0_register_file_0_n_112_283),.ZN(execution_unit_0_register_file_0_n_112_284));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_299 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[14]),.ZN(execution_unit_0_register_file_0_n_112_285));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_300 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[14]),.ZN(execution_unit_0_register_file_0_n_112_286));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_301 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[14]),.ZN(execution_unit_0_register_file_0_n_112_287));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_302 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[14]),.ZN(execution_unit_0_register_file_0_n_112_288));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_303 (.A1(execution_unit_0_register_file_0_n_112_285),.A2(execution_unit_0_register_file_0_n_112_286),.A3(execution_unit_0_register_file_0_n_112_287),.A4(execution_unit_0_register_file_0_n_112_288),.ZN(execution_unit_0_register_file_0_n_112_289));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_304 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[14]),.ZN(execution_unit_0_register_file_0_n_112_290));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_305 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[14]),.ZN(execution_unit_0_register_file_0_n_112_291));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_306 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[14]),.ZN(execution_unit_0_register_file_0_n_112_292));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_307 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[14]),.ZN(execution_unit_0_register_file_0_n_112_293));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_308 (.A1(execution_unit_0_register_file_0_n_112_290),.A2(execution_unit_0_register_file_0_n_112_291),.A3(execution_unit_0_register_file_0_n_112_292),.A4(execution_unit_0_register_file_0_n_112_293),.ZN(execution_unit_0_register_file_0_n_112_294));
	AND2_X1_LVT execution_unit_0register_file_0i_112_309 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[14]),.ZN(execution_unit_0_register_file_0_n_112_295));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_310 (.A1(execution_unit_0_register_file_0_n_112_284),.A2(execution_unit_0_register_file_0_n_112_289),.A3(execution_unit_0_register_file_0_n_112_294),.A4(execution_unit_0_register_file_0_n_112_295),.ZN(execution_unit_0_register_file_0_n_112_296));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_311 (.A1(inst_dest[0]),.A2(pc[14]),.ZN(execution_unit_0_register_file_0_n_112_297));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_312 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[14]),.ZN(execution_unit_0_register_file_0_n_112_298));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_313 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[14]),.ZN(execution_unit_0_register_file_0_n_112_299));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_314 (.A1(execution_unit_0_register_file_0_n_112_296),.A2(execution_unit_0_register_file_0_n_112_297),.A3(execution_unit_0_register_file_0_n_112_298),.A4(execution_unit_0_register_file_0_n_112_299),.ZN(dbg_reg_din[14]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_273 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[13]),.ZN(execution_unit_0_register_file_0_n_112_260));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_274 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[13]),.ZN(execution_unit_0_register_file_0_n_112_261));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_275 (.A1(inst_dest[2]),.A2(execution_unit_0_register_file_0_n_2),.ZN(execution_unit_0_register_file_0_n_112_262));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_276 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[13]),.ZN(execution_unit_0_register_file_0_n_112_263));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_277 (.A1(execution_unit_0_register_file_0_n_112_260),.A2(execution_unit_0_register_file_0_n_112_261),.A3(execution_unit_0_register_file_0_n_112_262),.A4(execution_unit_0_register_file_0_n_112_263),.ZN(execution_unit_0_register_file_0_n_112_264));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_278 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[13]),.ZN(execution_unit_0_register_file_0_n_112_265));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_279 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[13]),.ZN(execution_unit_0_register_file_0_n_112_266));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_280 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[13]),.ZN(execution_unit_0_register_file_0_n_112_267));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_281 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[13]),.ZN(execution_unit_0_register_file_0_n_112_268));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_282 (.A1(execution_unit_0_register_file_0_n_112_265),.A2(execution_unit_0_register_file_0_n_112_266),.A3(execution_unit_0_register_file_0_n_112_267),.A4(execution_unit_0_register_file_0_n_112_268),.ZN(execution_unit_0_register_file_0_n_112_269));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_283 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[13]),.ZN(execution_unit_0_register_file_0_n_112_270));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_284 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[13]),.ZN(execution_unit_0_register_file_0_n_112_271));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_285 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[13]),.ZN(execution_unit_0_register_file_0_n_112_272));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_286 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[13]),.ZN(execution_unit_0_register_file_0_n_112_273));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_287 (.A1(execution_unit_0_register_file_0_n_112_270),.A2(execution_unit_0_register_file_0_n_112_271),.A3(execution_unit_0_register_file_0_n_112_272),.A4(execution_unit_0_register_file_0_n_112_273),.ZN(execution_unit_0_register_file_0_n_112_274));
	AND2_X1_LVT execution_unit_0register_file_0i_112_288 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[13]),.ZN(execution_unit_0_register_file_0_n_112_275));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_289 (.A1(execution_unit_0_register_file_0_n_112_264),.A2(execution_unit_0_register_file_0_n_112_269),.A3(execution_unit_0_register_file_0_n_112_274),.A4(execution_unit_0_register_file_0_n_112_275),.ZN(execution_unit_0_register_file_0_n_112_276));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_290 (.A1(inst_dest[0]),.A2(pc[13]),.ZN(execution_unit_0_register_file_0_n_112_277));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_291 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[13]),.ZN(execution_unit_0_register_file_0_n_112_278));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_292 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[13]),.ZN(execution_unit_0_register_file_0_n_112_279));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_293 (.A1(execution_unit_0_register_file_0_n_112_276),.A2(execution_unit_0_register_file_0_n_112_277),.A3(execution_unit_0_register_file_0_n_112_278),.A4(execution_unit_0_register_file_0_n_112_279),.ZN(dbg_reg_din[13]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_252 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[12]),.ZN(execution_unit_0_register_file_0_n_112_240));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_253 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[12]),.ZN(execution_unit_0_register_file_0_n_112_241));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_254 (.A1(inst_dest[2]),.A2(execution_unit_0_register_file_0_n_3),.ZN(execution_unit_0_register_file_0_n_112_242));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_255 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[12]),.ZN(execution_unit_0_register_file_0_n_112_243));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_256 (.A1(execution_unit_0_register_file_0_n_112_240),.A2(execution_unit_0_register_file_0_n_112_241),.A3(execution_unit_0_register_file_0_n_112_242),.A4(execution_unit_0_register_file_0_n_112_243),.ZN(execution_unit_0_register_file_0_n_112_244));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_257 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[12]),.ZN(execution_unit_0_register_file_0_n_112_245));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_258 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[12]),.ZN(execution_unit_0_register_file_0_n_112_246));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_259 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[12]),.ZN(execution_unit_0_register_file_0_n_112_247));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_260 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[12]),.ZN(execution_unit_0_register_file_0_n_112_248));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_261 (.A1(execution_unit_0_register_file_0_n_112_245),.A2(execution_unit_0_register_file_0_n_112_246),.A3(execution_unit_0_register_file_0_n_112_247),.A4(execution_unit_0_register_file_0_n_112_248),.ZN(execution_unit_0_register_file_0_n_112_249));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_262 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[12]),.ZN(execution_unit_0_register_file_0_n_112_250));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_263 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[12]),.ZN(execution_unit_0_register_file_0_n_112_251));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_264 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[12]),.ZN(execution_unit_0_register_file_0_n_112_252));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_265 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[12]),.ZN(execution_unit_0_register_file_0_n_112_253));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_266 (.A1(execution_unit_0_register_file_0_n_112_250),.A2(execution_unit_0_register_file_0_n_112_251),.A3(execution_unit_0_register_file_0_n_112_252),.A4(execution_unit_0_register_file_0_n_112_253),.ZN(execution_unit_0_register_file_0_n_112_254));
	AND2_X1_LVT execution_unit_0register_file_0i_112_267 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[12]),.ZN(execution_unit_0_register_file_0_n_112_255));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_268 (.A1(execution_unit_0_register_file_0_n_112_244),.A2(execution_unit_0_register_file_0_n_112_249),.A3(execution_unit_0_register_file_0_n_112_254),.A4(execution_unit_0_register_file_0_n_112_255),.ZN(execution_unit_0_register_file_0_n_112_256));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_269 (.A1(inst_dest[0]),.A2(pc[12]),.ZN(execution_unit_0_register_file_0_n_112_257));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_270 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[12]),.ZN(execution_unit_0_register_file_0_n_112_258));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_271 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[12]),.ZN(execution_unit_0_register_file_0_n_112_259));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_272 (.A1(execution_unit_0_register_file_0_n_112_256),.A2(execution_unit_0_register_file_0_n_112_257),.A3(execution_unit_0_register_file_0_n_112_258),.A4(execution_unit_0_register_file_0_n_112_259),.ZN(dbg_reg_din[12]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_231 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[11]),.ZN(execution_unit_0_register_file_0_n_112_220));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_232 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[11]),.ZN(execution_unit_0_register_file_0_n_112_221));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_233 (.A1(inst_dest[2]),.A2(execution_unit_0_register_file_0_n_4),.ZN(execution_unit_0_register_file_0_n_112_222));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_234 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[11]),.ZN(execution_unit_0_register_file_0_n_112_223));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_235 (.A1(execution_unit_0_register_file_0_n_112_220),.A2(execution_unit_0_register_file_0_n_112_221),.A3(execution_unit_0_register_file_0_n_112_222),.A4(execution_unit_0_register_file_0_n_112_223),.ZN(execution_unit_0_register_file_0_n_112_224));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_236 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[11]),.ZN(execution_unit_0_register_file_0_n_112_225));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_237 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[11]),.ZN(execution_unit_0_register_file_0_n_112_226));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_238 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[11]),.ZN(execution_unit_0_register_file_0_n_112_227));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_239 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[11]),.ZN(execution_unit_0_register_file_0_n_112_228));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_240 (.A1(execution_unit_0_register_file_0_n_112_225),.A2(execution_unit_0_register_file_0_n_112_226),.A3(execution_unit_0_register_file_0_n_112_227),.A4(execution_unit_0_register_file_0_n_112_228),.ZN(execution_unit_0_register_file_0_n_112_229));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_241 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[11]),.ZN(execution_unit_0_register_file_0_n_112_230));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_242 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[11]),.ZN(execution_unit_0_register_file_0_n_112_231));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_243 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[11]),.ZN(execution_unit_0_register_file_0_n_112_232));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_244 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[11]),.ZN(execution_unit_0_register_file_0_n_112_233));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_245 (.A1(execution_unit_0_register_file_0_n_112_230),.A2(execution_unit_0_register_file_0_n_112_231),.A3(execution_unit_0_register_file_0_n_112_232),.A4(execution_unit_0_register_file_0_n_112_233),.ZN(execution_unit_0_register_file_0_n_112_234));
	AND2_X1_LVT execution_unit_0register_file_0i_112_246 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[11]),.ZN(execution_unit_0_register_file_0_n_112_235));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_247 (.A1(execution_unit_0_register_file_0_n_112_224),.A2(execution_unit_0_register_file_0_n_112_229),.A3(execution_unit_0_register_file_0_n_112_234),.A4(execution_unit_0_register_file_0_n_112_235),.ZN(execution_unit_0_register_file_0_n_112_236));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_248 (.A1(inst_dest[0]),.A2(pc[11]),.ZN(execution_unit_0_register_file_0_n_112_237));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_249 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[11]),.ZN(execution_unit_0_register_file_0_n_112_238));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_250 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[11]),.ZN(execution_unit_0_register_file_0_n_112_239));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_251 (.A1(execution_unit_0_register_file_0_n_112_236),.A2(execution_unit_0_register_file_0_n_112_237),.A3(execution_unit_0_register_file_0_n_112_238),.A4(execution_unit_0_register_file_0_n_112_239),.ZN(dbg_reg_din[11]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_210 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[10]),.ZN(execution_unit_0_register_file_0_n_112_200));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_211 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[10]),.ZN(execution_unit_0_register_file_0_n_112_201));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_212 (.A1(inst_dest[2]),.A2(execution_unit_0_register_file_0_n_5),.ZN(execution_unit_0_register_file_0_n_112_202));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_213 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[10]),.ZN(execution_unit_0_register_file_0_n_112_203));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_214 (.A1(execution_unit_0_register_file_0_n_112_200),.A2(execution_unit_0_register_file_0_n_112_201),.A3(execution_unit_0_register_file_0_n_112_202),.A4(execution_unit_0_register_file_0_n_112_203),.ZN(execution_unit_0_register_file_0_n_112_204));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_215 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[10]),.ZN(execution_unit_0_register_file_0_n_112_205));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_216 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[10]),.ZN(execution_unit_0_register_file_0_n_112_206));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_217 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[10]),.ZN(execution_unit_0_register_file_0_n_112_207));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_218 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[10]),.ZN(execution_unit_0_register_file_0_n_112_208));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_219 (.A1(execution_unit_0_register_file_0_n_112_205),.A2(execution_unit_0_register_file_0_n_112_206),.A3(execution_unit_0_register_file_0_n_112_207),.A4(execution_unit_0_register_file_0_n_112_208),.ZN(execution_unit_0_register_file_0_n_112_209));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_220 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[10]),.ZN(execution_unit_0_register_file_0_n_112_210));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_221 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[10]),.ZN(execution_unit_0_register_file_0_n_112_211));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_222 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[10]),.ZN(execution_unit_0_register_file_0_n_112_212));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_223 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[10]),.ZN(execution_unit_0_register_file_0_n_112_213));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_224 (.A1(execution_unit_0_register_file_0_n_112_210),.A2(execution_unit_0_register_file_0_n_112_211),.A3(execution_unit_0_register_file_0_n_112_212),.A4(execution_unit_0_register_file_0_n_112_213),.ZN(execution_unit_0_register_file_0_n_112_214));
	AND2_X1_LVT execution_unit_0register_file_0i_112_225 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[10]),.ZN(execution_unit_0_register_file_0_n_112_215));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_226 (.A1(execution_unit_0_register_file_0_n_112_204),.A2(execution_unit_0_register_file_0_n_112_209),.A3(execution_unit_0_register_file_0_n_112_214),.A4(execution_unit_0_register_file_0_n_112_215),.ZN(execution_unit_0_register_file_0_n_112_216));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_227 (.A1(inst_dest[0]),.A2(pc[10]),.ZN(execution_unit_0_register_file_0_n_112_217));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_228 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[10]),.ZN(execution_unit_0_register_file_0_n_112_218));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_229 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[10]),.ZN(execution_unit_0_register_file_0_n_112_219));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_230 (.A1(execution_unit_0_register_file_0_n_112_216),.A2(execution_unit_0_register_file_0_n_112_217),.A3(execution_unit_0_register_file_0_n_112_218),.A4(execution_unit_0_register_file_0_n_112_219),.ZN(dbg_reg_din[10]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_189 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[9]),.ZN(execution_unit_0_register_file_0_n_112_180));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_190 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[9]),.ZN(execution_unit_0_register_file_0_n_112_181));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_191 (.A1(inst_dest[2]),.A2(execution_unit_0_register_file_0_n_6),.ZN(execution_unit_0_register_file_0_n_112_182));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_192 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[9]),.ZN(execution_unit_0_register_file_0_n_112_183));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_193 (.A1(execution_unit_0_register_file_0_n_112_180),.A2(execution_unit_0_register_file_0_n_112_181),.A3(execution_unit_0_register_file_0_n_112_182),.A4(execution_unit_0_register_file_0_n_112_183),.ZN(execution_unit_0_register_file_0_n_112_184));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_194 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[9]),.ZN(execution_unit_0_register_file_0_n_112_185));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_195 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[9]),.ZN(execution_unit_0_register_file_0_n_112_186));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_196 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[9]),.ZN(execution_unit_0_register_file_0_n_112_187));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_197 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[9]),.ZN(execution_unit_0_register_file_0_n_112_188));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_198 (.A1(execution_unit_0_register_file_0_n_112_185),.A2(execution_unit_0_register_file_0_n_112_186),.A3(execution_unit_0_register_file_0_n_112_187),.A4(execution_unit_0_register_file_0_n_112_188),.ZN(execution_unit_0_register_file_0_n_112_189));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_199 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[9]),.ZN(execution_unit_0_register_file_0_n_112_190));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_200 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[9]),.ZN(execution_unit_0_register_file_0_n_112_191));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_201 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[9]),.ZN(execution_unit_0_register_file_0_n_112_192));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_202 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[9]),.ZN(execution_unit_0_register_file_0_n_112_193));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_203 (.A1(execution_unit_0_register_file_0_n_112_190),.A2(execution_unit_0_register_file_0_n_112_191),.A3(execution_unit_0_register_file_0_n_112_192),.A4(execution_unit_0_register_file_0_n_112_193),.ZN(execution_unit_0_register_file_0_n_112_194));
	AND2_X1_LVT execution_unit_0register_file_0i_112_204 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[9]),.ZN(execution_unit_0_register_file_0_n_112_195));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_205 (.A1(execution_unit_0_register_file_0_n_112_184),.A2(execution_unit_0_register_file_0_n_112_189),.A3(execution_unit_0_register_file_0_n_112_194),.A4(execution_unit_0_register_file_0_n_112_195),.ZN(execution_unit_0_register_file_0_n_112_196));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_206 (.A1(inst_dest[0]),.A2(pc[9]),.ZN(execution_unit_0_register_file_0_n_112_197));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_207 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[9]),.ZN(execution_unit_0_register_file_0_n_112_198));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_208 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[9]),.ZN(execution_unit_0_register_file_0_n_112_199));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_209 (.A1(execution_unit_0_register_file_0_n_112_196),.A2(execution_unit_0_register_file_0_n_112_197),.A3(execution_unit_0_register_file_0_n_112_198),.A4(execution_unit_0_register_file_0_n_112_199),.ZN(dbg_reg_din[9]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_168 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[8]),.ZN(execution_unit_0_register_file_0_n_112_160));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_169 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[8]),.ZN(execution_unit_0_register_file_0_n_112_161));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_170 (.A1(inst_dest[2]),.A2(execution_unit_0_status[3]),.ZN(execution_unit_0_register_file_0_n_112_162));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_171 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[8]),.ZN(execution_unit_0_register_file_0_n_112_163));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_172 (.A1(execution_unit_0_register_file_0_n_112_160),.A2(execution_unit_0_register_file_0_n_112_161),.A3(execution_unit_0_register_file_0_n_112_162),.A4(execution_unit_0_register_file_0_n_112_163),.ZN(execution_unit_0_register_file_0_n_112_164));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_173 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[8]),.ZN(execution_unit_0_register_file_0_n_112_165));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_174 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[8]),.ZN(execution_unit_0_register_file_0_n_112_166));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_175 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[8]),.ZN(execution_unit_0_register_file_0_n_112_167));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_176 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[8]),.ZN(execution_unit_0_register_file_0_n_112_168));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_177 (.A1(execution_unit_0_register_file_0_n_112_165),.A2(execution_unit_0_register_file_0_n_112_166),.A3(execution_unit_0_register_file_0_n_112_167),.A4(execution_unit_0_register_file_0_n_112_168),.ZN(execution_unit_0_register_file_0_n_112_169));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_178 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[8]),.ZN(execution_unit_0_register_file_0_n_112_170));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_179 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[8]),.ZN(execution_unit_0_register_file_0_n_112_171));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_180 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[8]),.ZN(execution_unit_0_register_file_0_n_112_172));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_181 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[8]),.ZN(execution_unit_0_register_file_0_n_112_173));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_182 (.A1(execution_unit_0_register_file_0_n_112_170),.A2(execution_unit_0_register_file_0_n_112_171),.A3(execution_unit_0_register_file_0_n_112_172),.A4(execution_unit_0_register_file_0_n_112_173),.ZN(execution_unit_0_register_file_0_n_112_174));
	AND2_X1_LVT execution_unit_0register_file_0i_112_183 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[8]),.ZN(execution_unit_0_register_file_0_n_112_175));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_184 (.A1(execution_unit_0_register_file_0_n_112_164),.A2(execution_unit_0_register_file_0_n_112_169),.A3(execution_unit_0_register_file_0_n_112_174),.A4(execution_unit_0_register_file_0_n_112_175),.ZN(execution_unit_0_register_file_0_n_112_176));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_185 (.A1(inst_dest[0]),.A2(pc[8]),.ZN(execution_unit_0_register_file_0_n_112_177));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_186 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[8]),.ZN(execution_unit_0_register_file_0_n_112_178));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_187 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[8]),.ZN(execution_unit_0_register_file_0_n_112_179));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_188 (.A1(execution_unit_0_register_file_0_n_112_176),.A2(execution_unit_0_register_file_0_n_112_177),.A3(execution_unit_0_register_file_0_n_112_178),.A4(execution_unit_0_register_file_0_n_112_179),.ZN(dbg_reg_din[8]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_147 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[7]),.ZN(execution_unit_0_register_file_0_n_112_140));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_148 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[7]),.ZN(execution_unit_0_register_file_0_n_112_141));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_149 (.A1(inst_dest[2]),.A2(scg1),.ZN(execution_unit_0_register_file_0_n_112_142));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_150 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[7]),.ZN(execution_unit_0_register_file_0_n_112_143));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_151 (.A1(execution_unit_0_register_file_0_n_112_140),.A2(execution_unit_0_register_file_0_n_112_141),.A3(execution_unit_0_register_file_0_n_112_142),.A4(execution_unit_0_register_file_0_n_112_143),.ZN(execution_unit_0_register_file_0_n_112_144));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_152 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[7]),.ZN(execution_unit_0_register_file_0_n_112_145));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_153 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[7]),.ZN(execution_unit_0_register_file_0_n_112_146));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_154 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[7]),.ZN(execution_unit_0_register_file_0_n_112_147));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_155 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[7]),.ZN(execution_unit_0_register_file_0_n_112_148));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_156 (.A1(execution_unit_0_register_file_0_n_112_145),.A2(execution_unit_0_register_file_0_n_112_146),.A3(execution_unit_0_register_file_0_n_112_147),.A4(execution_unit_0_register_file_0_n_112_148),.ZN(execution_unit_0_register_file_0_n_112_149));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_157 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[7]),.ZN(execution_unit_0_register_file_0_n_112_150));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_158 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[7]),.ZN(execution_unit_0_register_file_0_n_112_151));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_159 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[7]),.ZN(execution_unit_0_register_file_0_n_112_152));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_160 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[7]),.ZN(execution_unit_0_register_file_0_n_112_153));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_161 (.A1(execution_unit_0_register_file_0_n_112_150),.A2(execution_unit_0_register_file_0_n_112_151),.A3(execution_unit_0_register_file_0_n_112_152),.A4(execution_unit_0_register_file_0_n_112_153),.ZN(execution_unit_0_register_file_0_n_112_154));
	AND2_X1_LVT execution_unit_0register_file_0i_112_162 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[7]),.ZN(execution_unit_0_register_file_0_n_112_155));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_163 (.A1(execution_unit_0_register_file_0_n_112_144),.A2(execution_unit_0_register_file_0_n_112_149),.A3(execution_unit_0_register_file_0_n_112_154),.A4(execution_unit_0_register_file_0_n_112_155),.ZN(execution_unit_0_register_file_0_n_112_156));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_164 (.A1(inst_dest[0]),.A2(pc[7]),.ZN(execution_unit_0_register_file_0_n_112_157));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_165 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[7]),.ZN(execution_unit_0_register_file_0_n_112_158));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_166 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[7]),.ZN(execution_unit_0_register_file_0_n_112_159));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_167 (.A1(execution_unit_0_register_file_0_n_112_156),.A2(execution_unit_0_register_file_0_n_112_157),.A3(execution_unit_0_register_file_0_n_112_158),.A4(execution_unit_0_register_file_0_n_112_159),.ZN(dbg_reg_din[7]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_126 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[6]),.ZN(execution_unit_0_register_file_0_n_112_120));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_127 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[6]),.ZN(execution_unit_0_register_file_0_n_112_121));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_128 (.A1(inst_dest[2]),.A2(scg0),.ZN(execution_unit_0_register_file_0_n_112_122));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_129 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[6]),.ZN(execution_unit_0_register_file_0_n_112_123));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_130 (.A1(execution_unit_0_register_file_0_n_112_120),.A2(execution_unit_0_register_file_0_n_112_121),.A3(execution_unit_0_register_file_0_n_112_122),.A4(execution_unit_0_register_file_0_n_112_123),.ZN(execution_unit_0_register_file_0_n_112_124));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_131 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[6]),.ZN(execution_unit_0_register_file_0_n_112_125));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_132 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[6]),.ZN(execution_unit_0_register_file_0_n_112_126));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_133 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[6]),.ZN(execution_unit_0_register_file_0_n_112_127));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_134 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[6]),.ZN(execution_unit_0_register_file_0_n_112_128));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_135 (.A1(execution_unit_0_register_file_0_n_112_125),.A2(execution_unit_0_register_file_0_n_112_126),.A3(execution_unit_0_register_file_0_n_112_127),.A4(execution_unit_0_register_file_0_n_112_128),.ZN(execution_unit_0_register_file_0_n_112_129));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_136 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[6]),.ZN(execution_unit_0_register_file_0_n_112_130));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_137 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[6]),.ZN(execution_unit_0_register_file_0_n_112_131));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_138 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[6]),.ZN(execution_unit_0_register_file_0_n_112_132));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_139 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[6]),.ZN(execution_unit_0_register_file_0_n_112_133));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_140 (.A1(execution_unit_0_register_file_0_n_112_130),.A2(execution_unit_0_register_file_0_n_112_131),.A3(execution_unit_0_register_file_0_n_112_132),.A4(execution_unit_0_register_file_0_n_112_133),.ZN(execution_unit_0_register_file_0_n_112_134));
	AND2_X1_LVT execution_unit_0register_file_0i_112_141 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[6]),.ZN(execution_unit_0_register_file_0_n_112_135));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_142 (.A1(execution_unit_0_register_file_0_n_112_124),.A2(execution_unit_0_register_file_0_n_112_129),.A3(execution_unit_0_register_file_0_n_112_134),.A4(execution_unit_0_register_file_0_n_112_135),.ZN(execution_unit_0_register_file_0_n_112_136));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_143 (.A1(inst_dest[0]),.A2(pc[6]),.ZN(execution_unit_0_register_file_0_n_112_137));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_144 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[6]),.ZN(execution_unit_0_register_file_0_n_112_138));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_145 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[6]),.ZN(execution_unit_0_register_file_0_n_112_139));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_146 (.A1(execution_unit_0_register_file_0_n_112_136),.A2(execution_unit_0_register_file_0_n_112_137),.A3(execution_unit_0_register_file_0_n_112_138),.A4(execution_unit_0_register_file_0_n_112_139),.ZN(dbg_reg_din[6]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_105 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[5]),.ZN(execution_unit_0_register_file_0_n_112_100));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_106 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[5]),.ZN(execution_unit_0_register_file_0_n_112_101));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_107 (.A1(inst_dest[2]),.A2(oscoff),.ZN(execution_unit_0_register_file_0_n_112_102));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_108 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[5]),.ZN(execution_unit_0_register_file_0_n_112_103));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_109 (.A1(execution_unit_0_register_file_0_n_112_100),.A2(execution_unit_0_register_file_0_n_112_101),.A3(execution_unit_0_register_file_0_n_112_102),.A4(execution_unit_0_register_file_0_n_112_103),.ZN(execution_unit_0_register_file_0_n_112_104));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_110 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[5]),.ZN(execution_unit_0_register_file_0_n_112_105));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_111 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[5]),.ZN(execution_unit_0_register_file_0_n_112_106));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_112 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[5]),.ZN(execution_unit_0_register_file_0_n_112_107));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_113 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[5]),.ZN(execution_unit_0_register_file_0_n_112_108));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_114 (.A1(execution_unit_0_register_file_0_n_112_105),.A2(execution_unit_0_register_file_0_n_112_106),.A3(execution_unit_0_register_file_0_n_112_107),.A4(execution_unit_0_register_file_0_n_112_108),.ZN(execution_unit_0_register_file_0_n_112_109));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_115 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[5]),.ZN(execution_unit_0_register_file_0_n_112_110));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_116 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[5]),.ZN(execution_unit_0_register_file_0_n_112_111));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_117 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[5]),.ZN(execution_unit_0_register_file_0_n_112_112));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_118 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[5]),.ZN(execution_unit_0_register_file_0_n_112_113));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_119 (.A1(execution_unit_0_register_file_0_n_112_110),.A2(execution_unit_0_register_file_0_n_112_111),.A3(execution_unit_0_register_file_0_n_112_112),.A4(execution_unit_0_register_file_0_n_112_113),.ZN(execution_unit_0_register_file_0_n_112_114));
	AND2_X1_LVT execution_unit_0register_file_0i_112_120 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[5]),.ZN(execution_unit_0_register_file_0_n_112_115));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_121 (.A1(execution_unit_0_register_file_0_n_112_104),.A2(execution_unit_0_register_file_0_n_112_109),.A3(execution_unit_0_register_file_0_n_112_114),.A4(execution_unit_0_register_file_0_n_112_115),.ZN(execution_unit_0_register_file_0_n_112_116));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_122 (.A1(inst_dest[0]),.A2(pc[5]),.ZN(execution_unit_0_register_file_0_n_112_117));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_123 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[5]),.ZN(execution_unit_0_register_file_0_n_112_118));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_124 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[5]),.ZN(execution_unit_0_register_file_0_n_112_119));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_125 (.A1(execution_unit_0_register_file_0_n_112_116),.A2(execution_unit_0_register_file_0_n_112_117),.A3(execution_unit_0_register_file_0_n_112_118),.A4(execution_unit_0_register_file_0_n_112_119),.ZN(dbg_reg_din[5]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_84 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[4]),.ZN(execution_unit_0_register_file_0_n_112_80));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_85 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[4]),.ZN(execution_unit_0_register_file_0_n_112_81));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_86 (.A1(inst_dest[2]),.A2(execution_unit_0_register_file_0_n_7),.ZN(execution_unit_0_register_file_0_n_112_82));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_87 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[4]),.ZN(execution_unit_0_register_file_0_n_112_83));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_88 (.A1(execution_unit_0_register_file_0_n_112_80),.A2(execution_unit_0_register_file_0_n_112_81),.A3(execution_unit_0_register_file_0_n_112_82),.A4(execution_unit_0_register_file_0_n_112_83),.ZN(execution_unit_0_register_file_0_n_112_84));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_89 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[4]),.ZN(execution_unit_0_register_file_0_n_112_85));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_90 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[4]),.ZN(execution_unit_0_register_file_0_n_112_86));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_91 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[4]),.ZN(execution_unit_0_register_file_0_n_112_87));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_92 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[4]),.ZN(execution_unit_0_register_file_0_n_112_88));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_93 (.A1(execution_unit_0_register_file_0_n_112_85),.A2(execution_unit_0_register_file_0_n_112_86),.A3(execution_unit_0_register_file_0_n_112_87),.A4(execution_unit_0_register_file_0_n_112_88),.ZN(execution_unit_0_register_file_0_n_112_89));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_94 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[4]),.ZN(execution_unit_0_register_file_0_n_112_90));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_95 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[4]),.ZN(execution_unit_0_register_file_0_n_112_91));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_96 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[4]),.ZN(execution_unit_0_register_file_0_n_112_92));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_97 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[4]),.ZN(execution_unit_0_register_file_0_n_112_93));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_98 (.A1(execution_unit_0_register_file_0_n_112_90),.A2(execution_unit_0_register_file_0_n_112_91),.A3(execution_unit_0_register_file_0_n_112_92),.A4(execution_unit_0_register_file_0_n_112_93),.ZN(execution_unit_0_register_file_0_n_112_94));
	AND2_X1_LVT execution_unit_0register_file_0i_112_99 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[4]),.ZN(execution_unit_0_register_file_0_n_112_95));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_100 (.A1(execution_unit_0_register_file_0_n_112_84),.A2(execution_unit_0_register_file_0_n_112_89),.A3(execution_unit_0_register_file_0_n_112_94),.A4(execution_unit_0_register_file_0_n_112_95),.ZN(execution_unit_0_register_file_0_n_112_96));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_101 (.A1(inst_dest[0]),.A2(pc[4]),.ZN(execution_unit_0_register_file_0_n_112_97));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_102 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[4]),.ZN(execution_unit_0_register_file_0_n_112_98));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_103 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[4]),.ZN(execution_unit_0_register_file_0_n_112_99));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_104 (.A1(execution_unit_0_register_file_0_n_112_96),.A2(execution_unit_0_register_file_0_n_112_97),.A3(execution_unit_0_register_file_0_n_112_98),.A4(execution_unit_0_register_file_0_n_112_99),.ZN(dbg_reg_din[4]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_63 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[3]),.ZN(execution_unit_0_register_file_0_n_112_60));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_64 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[3]),.ZN(execution_unit_0_register_file_0_n_112_61));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_65 (.A1(inst_dest[2]),.A2(gie),.ZN(execution_unit_0_register_file_0_n_112_62));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_66 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[3]),.ZN(execution_unit_0_register_file_0_n_112_63));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_67 (.A1(execution_unit_0_register_file_0_n_112_60),.A2(execution_unit_0_register_file_0_n_112_61),.A3(execution_unit_0_register_file_0_n_112_62),.A4(execution_unit_0_register_file_0_n_112_63),.ZN(execution_unit_0_register_file_0_n_112_64));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_68 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[3]),.ZN(execution_unit_0_register_file_0_n_112_65));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_69 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[3]),.ZN(execution_unit_0_register_file_0_n_112_66));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_70 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[3]),.ZN(execution_unit_0_register_file_0_n_112_67));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_71 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[3]),.ZN(execution_unit_0_register_file_0_n_112_68));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_72 (.A1(execution_unit_0_register_file_0_n_112_65),.A2(execution_unit_0_register_file_0_n_112_66),.A3(execution_unit_0_register_file_0_n_112_67),.A4(execution_unit_0_register_file_0_n_112_68),.ZN(execution_unit_0_register_file_0_n_112_69));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_73 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[3]),.ZN(execution_unit_0_register_file_0_n_112_70));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_74 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[3]),.ZN(execution_unit_0_register_file_0_n_112_71));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_75 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[3]),.ZN(execution_unit_0_register_file_0_n_112_72));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_76 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[3]),.ZN(execution_unit_0_register_file_0_n_112_73));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_77 (.A1(execution_unit_0_register_file_0_n_112_70),.A2(execution_unit_0_register_file_0_n_112_71),.A3(execution_unit_0_register_file_0_n_112_72),.A4(execution_unit_0_register_file_0_n_112_73),.ZN(execution_unit_0_register_file_0_n_112_74));
	AND2_X1_LVT execution_unit_0register_file_0i_112_78 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[3]),.ZN(execution_unit_0_register_file_0_n_112_75));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_79 (.A1(execution_unit_0_register_file_0_n_112_64),.A2(execution_unit_0_register_file_0_n_112_69),.A3(execution_unit_0_register_file_0_n_112_74),.A4(execution_unit_0_register_file_0_n_112_75),.ZN(execution_unit_0_register_file_0_n_112_76));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_80 (.A1(inst_dest[0]),.A2(pc[3]),.ZN(execution_unit_0_register_file_0_n_112_77));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_81 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[3]),.ZN(execution_unit_0_register_file_0_n_112_78));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_82 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[3]),.ZN(execution_unit_0_register_file_0_n_112_79));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_83 (.A1(execution_unit_0_register_file_0_n_112_76),.A2(execution_unit_0_register_file_0_n_112_77),.A3(execution_unit_0_register_file_0_n_112_78),.A4(execution_unit_0_register_file_0_n_112_79),.ZN(dbg_reg_din[3]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_42 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[2]),.ZN(execution_unit_0_register_file_0_n_112_40));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_43 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[2]),.ZN(execution_unit_0_register_file_0_n_112_41));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_44 (.A1(inst_dest[2]),.A2(execution_unit_0_status[2]),.ZN(execution_unit_0_register_file_0_n_112_42));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_45 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[2]),.ZN(execution_unit_0_register_file_0_n_112_43));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_46 (.A1(execution_unit_0_register_file_0_n_112_40),.A2(execution_unit_0_register_file_0_n_112_41),.A3(execution_unit_0_register_file_0_n_112_42),.A4(execution_unit_0_register_file_0_n_112_43),.ZN(execution_unit_0_register_file_0_n_112_44));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_47 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[2]),.ZN(execution_unit_0_register_file_0_n_112_45));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_48 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[2]),.ZN(execution_unit_0_register_file_0_n_112_46));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_49 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[2]),.ZN(execution_unit_0_register_file_0_n_112_47));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_50 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[2]),.ZN(execution_unit_0_register_file_0_n_112_48));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_51 (.A1(execution_unit_0_register_file_0_n_112_45),.A2(execution_unit_0_register_file_0_n_112_46),.A3(execution_unit_0_register_file_0_n_112_47),.A4(execution_unit_0_register_file_0_n_112_48),.ZN(execution_unit_0_register_file_0_n_112_49));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_52 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[2]),.ZN(execution_unit_0_register_file_0_n_112_50));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_53 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[2]),.ZN(execution_unit_0_register_file_0_n_112_51));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_54 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[2]),.ZN(execution_unit_0_register_file_0_n_112_52));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_55 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[2]),.ZN(execution_unit_0_register_file_0_n_112_53));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_56 (.A1(execution_unit_0_register_file_0_n_112_50),.A2(execution_unit_0_register_file_0_n_112_51),.A3(execution_unit_0_register_file_0_n_112_52),.A4(execution_unit_0_register_file_0_n_112_53),.ZN(execution_unit_0_register_file_0_n_112_54));
	AND2_X1_LVT execution_unit_0register_file_0i_112_57 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[2]),.ZN(execution_unit_0_register_file_0_n_112_55));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_58 (.A1(execution_unit_0_register_file_0_n_112_44),.A2(execution_unit_0_register_file_0_n_112_49),.A3(execution_unit_0_register_file_0_n_112_54),.A4(execution_unit_0_register_file_0_n_112_55),.ZN(execution_unit_0_register_file_0_n_112_56));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_59 (.A1(inst_dest[0]),.A2(pc[2]),.ZN(execution_unit_0_register_file_0_n_112_57));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_60 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[2]),.ZN(execution_unit_0_register_file_0_n_112_58));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_61 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[2]),.ZN(execution_unit_0_register_file_0_n_112_59));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_62 (.A1(execution_unit_0_register_file_0_n_112_56),.A2(execution_unit_0_register_file_0_n_112_57),.A3(execution_unit_0_register_file_0_n_112_58),.A4(execution_unit_0_register_file_0_n_112_59),.ZN(dbg_reg_din[2]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_21 (.A1(inst_dest[4]),.A2(execution_unit_0_register_file_0_r4[1]),.ZN(execution_unit_0_register_file_0_n_112_20));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_22 (.A1(inst_dest[3]),.A2(execution_unit_0_register_file_0_r3[1]),.ZN(execution_unit_0_register_file_0_n_112_21));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_23 (.A1(inst_dest[2]),.A2(execution_unit_0_status[1]),.ZN(execution_unit_0_register_file_0_n_112_22));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_24 (.A1(inst_dest[1]),.A2(execution_unit_0_register_file_0_r1[1]),.ZN(execution_unit_0_register_file_0_n_112_23));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_25 (.A1(execution_unit_0_register_file_0_n_112_20),.A2(execution_unit_0_register_file_0_n_112_21),.A3(execution_unit_0_register_file_0_n_112_22),.A4(execution_unit_0_register_file_0_n_112_23),.ZN(execution_unit_0_register_file_0_n_112_24));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_26 (.A1(inst_dest[12]),.A2(execution_unit_0_register_file_0_r12[1]),.ZN(execution_unit_0_register_file_0_n_112_25));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_27 (.A1(inst_dest[11]),.A2(execution_unit_0_register_file_0_r11[1]),.ZN(execution_unit_0_register_file_0_n_112_26));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_28 (.A1(inst_dest[10]),.A2(execution_unit_0_register_file_0_r10[1]),.ZN(execution_unit_0_register_file_0_n_112_27));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_29 (.A1(inst_dest[9]),.A2(execution_unit_0_register_file_0_r9[1]),.ZN(execution_unit_0_register_file_0_n_112_28));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_30 (.A1(execution_unit_0_register_file_0_n_112_25),.A2(execution_unit_0_register_file_0_n_112_26),.A3(execution_unit_0_register_file_0_n_112_27),.A4(execution_unit_0_register_file_0_n_112_28),.ZN(execution_unit_0_register_file_0_n_112_29));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_31 (.A1(inst_dest[8]),.A2(execution_unit_0_register_file_0_r8[1]),.ZN(execution_unit_0_register_file_0_n_112_30));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_32 (.A1(inst_dest[7]),.A2(execution_unit_0_register_file_0_r7[1]),.ZN(execution_unit_0_register_file_0_n_112_31));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_33 (.A1(inst_dest[6]),.A2(execution_unit_0_register_file_0_r6[1]),.ZN(execution_unit_0_register_file_0_n_112_32));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_34 (.A1(inst_dest[5]),.A2(execution_unit_0_register_file_0_r5[1]),.ZN(execution_unit_0_register_file_0_n_112_33));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_35 (.A1(execution_unit_0_register_file_0_n_112_30),.A2(execution_unit_0_register_file_0_n_112_31),.A3(execution_unit_0_register_file_0_n_112_32),.A4(execution_unit_0_register_file_0_n_112_33),.ZN(execution_unit_0_register_file_0_n_112_34));
	AND2_X1_LVT execution_unit_0register_file_0i_112_36 (.A1(inst_dest[13]),.A2(execution_unit_0_register_file_0_r13[1]),.ZN(execution_unit_0_register_file_0_n_112_35));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_37 (.A1(execution_unit_0_register_file_0_n_112_24),.A2(execution_unit_0_register_file_0_n_112_29),.A3(execution_unit_0_register_file_0_n_112_34),.A4(execution_unit_0_register_file_0_n_112_35),.ZN(execution_unit_0_register_file_0_n_112_36));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_38 (.A1(inst_dest[0]),.A2(pc[1]),.ZN(execution_unit_0_register_file_0_n_112_37));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_39 (.A1(inst_dest[15]),.A2(execution_unit_0_register_file_0_r15[1]),.ZN(execution_unit_0_register_file_0_n_112_38));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_40 (.A1(inst_dest[14]),.A2(execution_unit_0_register_file_0_r14[1]),.ZN(execution_unit_0_register_file_0_n_112_39));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_41 (.A1(execution_unit_0_register_file_0_n_112_36),.A2(execution_unit_0_register_file_0_n_112_37),.A3(execution_unit_0_register_file_0_n_112_38),.A4(execution_unit_0_register_file_0_n_112_39),.ZN(dbg_reg_din[1]));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_0 (.A1(execution_unit_0_register_file_0_r4[0]),.A2(inst_dest[4]),.ZN(execution_unit_0_register_file_0_n_112_0));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_1 (.A1(execution_unit_0_register_file_0_r3[0]),.A2(inst_dest[3]),.ZN(execution_unit_0_register_file_0_n_112_1));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_2 (.A1(execution_unit_0_status[0]),.A2(inst_dest[2]),.ZN(execution_unit_0_register_file_0_n_112_2));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_3 (.A1(execution_unit_0_register_file_0_r1[0]),.A2(inst_dest[1]),.ZN(execution_unit_0_register_file_0_n_112_3));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_4 (.A1(execution_unit_0_register_file_0_n_112_0),.A2(execution_unit_0_register_file_0_n_112_1),.A3(execution_unit_0_register_file_0_n_112_2),.A4(execution_unit_0_register_file_0_n_112_3),.ZN(execution_unit_0_register_file_0_n_112_4));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_5 (.A1(execution_unit_0_register_file_0_r12[0]),.A2(inst_dest[12]),.ZN(execution_unit_0_register_file_0_n_112_5));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_6 (.A1(execution_unit_0_register_file_0_r11[0]),.A2(inst_dest[11]),.ZN(execution_unit_0_register_file_0_n_112_6));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_7 (.A1(execution_unit_0_register_file_0_r10[0]),.A2(inst_dest[10]),.ZN(execution_unit_0_register_file_0_n_112_7));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_8 (.A1(execution_unit_0_register_file_0_r9[0]),.A2(inst_dest[9]),.ZN(execution_unit_0_register_file_0_n_112_8));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_9 (.A1(execution_unit_0_register_file_0_n_112_5),.A2(execution_unit_0_register_file_0_n_112_6),.A3(execution_unit_0_register_file_0_n_112_7),.A4(execution_unit_0_register_file_0_n_112_8),.ZN(execution_unit_0_register_file_0_n_112_9));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_10 (.A1(execution_unit_0_register_file_0_r8[0]),.A2(inst_dest[8]),.ZN(execution_unit_0_register_file_0_n_112_10));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_11 (.A1(execution_unit_0_register_file_0_r7[0]),.A2(inst_dest[7]),.ZN(execution_unit_0_register_file_0_n_112_11));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_12 (.A1(execution_unit_0_register_file_0_r6[0]),.A2(inst_dest[6]),.ZN(execution_unit_0_register_file_0_n_112_12));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_13 (.A1(execution_unit_0_register_file_0_r5[0]),.A2(inst_dest[5]),.ZN(execution_unit_0_register_file_0_n_112_13));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_14 (.A1(execution_unit_0_register_file_0_n_112_10),.A2(execution_unit_0_register_file_0_n_112_11),.A3(execution_unit_0_register_file_0_n_112_12),.A4(execution_unit_0_register_file_0_n_112_13),.ZN(execution_unit_0_register_file_0_n_112_14));
	AND2_X1_LVT execution_unit_0register_file_0i_112_15 (.A1(execution_unit_0_register_file_0_r13[0]),.A2(inst_dest[13]),.ZN(execution_unit_0_register_file_0_n_112_15));
	NOR4_X1_LVT execution_unit_0register_file_0i_112_16 (.A1(execution_unit_0_register_file_0_n_112_4),.A2(execution_unit_0_register_file_0_n_112_9),.A3(execution_unit_0_register_file_0_n_112_14),.A4(execution_unit_0_register_file_0_n_112_15),.ZN(execution_unit_0_register_file_0_n_112_16));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_17 (.A1(pc[0]),.A2(inst_dest[0]),.ZN(execution_unit_0_register_file_0_n_112_17));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_18 (.A1(execution_unit_0_register_file_0_r15[0]),.A2(inst_dest[15]),.ZN(execution_unit_0_register_file_0_n_112_18));
	NAND2_X1_LVT execution_unit_0register_file_0i_112_19 (.A1(execution_unit_0_register_file_0_r14[0]),.A2(inst_dest[14]),.ZN(execution_unit_0_register_file_0_n_112_19));
	NAND4_X1_LVT execution_unit_0register_file_0i_112_20 (.A1(execution_unit_0_register_file_0_n_112_16),.A2(execution_unit_0_register_file_0_n_112_17),.A3(execution_unit_0_register_file_0_n_112_18),.A4(execution_unit_0_register_file_0_n_112_19),.ZN(dbg_reg_din[0]));
	OR2_X1_LVT execution_unit_0i_8_0 (.A1(inst_bw),.A2(inst_alu[11]),.ZN(execution_unit_0_n_8_0));
	INV_X1_LVT execution_unit_0i_8_1 (.A(inst_alu[11]),.ZN(execution_unit_0_n_8_1));
	NAND2_X1_LVT execution_unit_0i_8_2 (.A1(execution_unit_0_n_8_1),.A2(inst_bw),.ZN(execution_unit_0_n_8_2));
	INV_X1_LVT execution_unit_0i_8_4 (.A(eu_mab[0]),.ZN(execution_unit_0_n_8_3));
	OAI21_X1_LVT execution_unit_0i_8_5 (.A(execution_unit_0_n_8_0),.B1(execution_unit_0_n_8_2),.B2(execution_unit_0_n_8_3),.ZN(execution_unit_0_n_15));
	AND2_X1_LVT execution_unit_0i_9_1 (.A1(execution_unit_0_mb_wr_det),.A2(execution_unit_0_n_15),.ZN(eu_mb_wr[1]));
	OAI21_X1_LVT execution_unit_0i_8_3 (.A(execution_unit_0_n_8_0),.B1(execution_unit_0_n_8_2),.B2(eu_mab[0]),.ZN(execution_unit_0_n_14));
	AND2_X1_LVT execution_unit_0i_9_0 (.A1(execution_unit_0_mb_wr_det),.A2(execution_unit_0_n_14),.ZN(eu_mb_wr[0]));
	INV_X1_LVT execution_unit_0i_17_0 (.A(inst_bw),.ZN(execution_unit_0_n_17_0));
	NAND2_X1_LVT execution_unit_0i_13_0 (.A1(e_state[0]),.A2(e_state[3]),.ZN(execution_unit_0_n_13_0));
	NOR3_X1_LVT execution_unit_0i_13_1 (.A1(execution_unit_0_n_13_0),.A2(e_state[1]),.A3(e_state[2]),.ZN(execution_unit_0_n_13_1));
	INV_X1_LVT execution_unit_0i_13_2 (.A(execution_unit_0_n_13_1),.ZN(execution_unit_0_n_13_2));
	AOI22_X1_LVT execution_unit_0i_13_33 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[15]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[15]),.ZN(execution_unit_0_n_13_18));
	INV_X1_LVT execution_unit_0i_13_34 (.A(execution_unit_0_n_13_18),.ZN(execution_unit_0_n_34));
	INV_X1_LVT execution_unit_0i_14_0 (.A(inst_so[5]),.ZN(execution_unit_0_n_14_0));
	AOI211_X1_LVT execution_unit_0i_14_1 (.A(execution_unit_0_n_7),.B(execution_unit_0_reg_sr_clr),.C1(execution_unit_0_n_14_0),.C2(execution_unit_0_n_0),.ZN(execution_unit_0_n_14_1));
	INV_X1_LVT execution_unit_0i_14_2 (.A(execution_unit_0_n_14_1),.ZN(execution_unit_0_n_35));
	INV_X1_LVT execution_unit_0i_15_3 (.A(execution_unit_0_n_35),.ZN(execution_unit_0_n_15_3));
	NAND2_X1_LVT execution_unit_0i_15_0 (.A1(e_state[0]),.A2(e_state[3]),.ZN(execution_unit_0_n_15_0));
	NOR3_X1_LVT execution_unit_0i_15_1 (.A1(execution_unit_0_n_15_0),.A2(e_state[1]),.A3(e_state[2]),.ZN(execution_unit_0_n_15_1));
	INV_X1_LVT execution_unit_0i_15_2 (.A(execution_unit_0_n_15_1),.ZN(execution_unit_0_n_15_2));
	NAND2_X1_LVT execution_unit_0i_15_4 (.A1(execution_unit_0_n_15_3),.A2(execution_unit_0_n_15_2),.ZN(execution_unit_0_n_36));
	CLKGATETST_X1_LVT execution_unit_0clk_gate_mdb_out_nxt_reg (.CK(cpu_mclk),.E(execution_unit_0_n_36),.SE(1'b0),.GCK(execution_unit_0_n_17));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b15___05F05d (.D(execution_unit_0_n_34),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(execution_unit_0_mdb_out_nxt[15]),.QN());
	AOI22_X1_LVT execution_unit_0i_13_17 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[7]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[7]),.ZN(execution_unit_0_n_13_10));
	INV_X1_LVT execution_unit_0i_13_18 (.A(execution_unit_0_n_13_10),.ZN(execution_unit_0_n_26));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b7___05F05d (.D(execution_unit_0_n_26),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(eu_mdb_out[7]),.QN());
	AOI22_X1_LVT execution_unit_0i_17_15 (.A1(execution_unit_0_n_17_0),.A2(execution_unit_0_mdb_out_nxt[15]),.B1(inst_bw),.B2(eu_mdb_out[7]),.ZN(execution_unit_0_n_17_8));
	INV_X1_LVT execution_unit_0i_17_16 (.A(execution_unit_0_n_17_8),.ZN(eu_mdb_out[15]));
	AOI22_X1_LVT execution_unit_0i_13_31 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[14]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[14]),.ZN(execution_unit_0_n_13_17));
	INV_X1_LVT execution_unit_0i_13_32 (.A(execution_unit_0_n_13_17),.ZN(execution_unit_0_n_33));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b14___05F05d (.D(execution_unit_0_n_33),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(execution_unit_0_mdb_out_nxt[14]),.QN());
	AOI22_X1_LVT execution_unit_0i_13_15 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[6]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[6]),.ZN(execution_unit_0_n_13_9));
	INV_X1_LVT execution_unit_0i_13_16 (.A(execution_unit_0_n_13_9),.ZN(execution_unit_0_n_25));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b6___05F05d (.D(execution_unit_0_n_25),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(eu_mdb_out[6]),.QN());
	AOI22_X1_LVT execution_unit_0i_17_13 (.A1(execution_unit_0_n_17_0),.A2(execution_unit_0_mdb_out_nxt[14]),.B1(inst_bw),.B2(eu_mdb_out[6]),.ZN(execution_unit_0_n_17_7));
	INV_X1_LVT execution_unit_0i_17_14 (.A(execution_unit_0_n_17_7),.ZN(eu_mdb_out[14]));
	AOI22_X1_LVT execution_unit_0i_13_29 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[13]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[13]),.ZN(execution_unit_0_n_13_16));
	INV_X1_LVT execution_unit_0i_13_30 (.A(execution_unit_0_n_13_16),.ZN(execution_unit_0_n_32));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b13___05F05d (.D(execution_unit_0_n_32),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(execution_unit_0_mdb_out_nxt[13]),.QN());
	AOI22_X1_LVT execution_unit_0i_13_13 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[5]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[5]),.ZN(execution_unit_0_n_13_8));
	INV_X1_LVT execution_unit_0i_13_14 (.A(execution_unit_0_n_13_8),.ZN(execution_unit_0_n_24));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b5___05F05d (.D(execution_unit_0_n_24),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(eu_mdb_out[5]),.QN());
	AOI22_X1_LVT execution_unit_0i_17_11 (.A1(execution_unit_0_n_17_0),.A2(execution_unit_0_mdb_out_nxt[13]),.B1(inst_bw),.B2(eu_mdb_out[5]),.ZN(execution_unit_0_n_17_6));
	INV_X1_LVT execution_unit_0i_17_12 (.A(execution_unit_0_n_17_6),.ZN(eu_mdb_out[13]));
	AOI22_X1_LVT execution_unit_0i_13_27 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[12]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[12]),.ZN(execution_unit_0_n_13_15));
	INV_X1_LVT execution_unit_0i_13_28 (.A(execution_unit_0_n_13_15),.ZN(execution_unit_0_n_31));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b12___05F05d (.D(execution_unit_0_n_31),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(execution_unit_0_mdb_out_nxt[12]),.QN());
	AOI22_X1_LVT execution_unit_0i_13_11 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[4]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[4]),.ZN(execution_unit_0_n_13_7));
	INV_X1_LVT execution_unit_0i_13_12 (.A(execution_unit_0_n_13_7),.ZN(execution_unit_0_n_23));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b4___05F05d (.D(execution_unit_0_n_23),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(eu_mdb_out[4]),.QN());
	AOI22_X1_LVT execution_unit_0i_17_9 (.A1(execution_unit_0_n_17_0),.A2(execution_unit_0_mdb_out_nxt[12]),.B1(inst_bw),.B2(eu_mdb_out[4]),.ZN(execution_unit_0_n_17_5));
	INV_X1_LVT execution_unit_0i_17_10 (.A(execution_unit_0_n_17_5),.ZN(eu_mdb_out[12]));
	AOI22_X1_LVT execution_unit_0i_13_25 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[11]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[11]),.ZN(execution_unit_0_n_13_14));
	INV_X1_LVT execution_unit_0i_13_26 (.A(execution_unit_0_n_13_14),.ZN(execution_unit_0_n_30));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b11___05F05d (.D(execution_unit_0_n_30),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(execution_unit_0_mdb_out_nxt[11]),.QN());
	AOI22_X1_LVT execution_unit_0i_13_9 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[3]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[3]),.ZN(execution_unit_0_n_13_6));
	INV_X1_LVT execution_unit_0i_13_10 (.A(execution_unit_0_n_13_6),.ZN(execution_unit_0_n_22));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b3___05F05d (.D(execution_unit_0_n_22),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(eu_mdb_out[3]),.QN());
	AOI22_X1_LVT execution_unit_0i_17_7 (.A1(execution_unit_0_n_17_0),.A2(execution_unit_0_mdb_out_nxt[11]),.B1(inst_bw),.B2(eu_mdb_out[3]),.ZN(execution_unit_0_n_17_4));
	INV_X1_LVT execution_unit_0i_17_8 (.A(execution_unit_0_n_17_4),.ZN(eu_mdb_out[11]));
	AOI22_X1_LVT execution_unit_0i_13_23 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[10]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[10]),.ZN(execution_unit_0_n_13_13));
	INV_X1_LVT execution_unit_0i_13_24 (.A(execution_unit_0_n_13_13),.ZN(execution_unit_0_n_29));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b10___05F05d (.D(execution_unit_0_n_29),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(execution_unit_0_mdb_out_nxt[10]),.QN());
	AOI22_X1_LVT execution_unit_0i_13_7 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[2]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[2]),.ZN(execution_unit_0_n_13_5));
	INV_X1_LVT execution_unit_0i_13_8 (.A(execution_unit_0_n_13_5),.ZN(execution_unit_0_n_21));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b2___05F05d (.D(execution_unit_0_n_21),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(eu_mdb_out[2]),.QN());
	AOI22_X1_LVT execution_unit_0i_17_5 (.A1(execution_unit_0_n_17_0),.A2(execution_unit_0_mdb_out_nxt[10]),.B1(inst_bw),.B2(eu_mdb_out[2]),.ZN(execution_unit_0_n_17_3));
	INV_X1_LVT execution_unit_0i_17_6 (.A(execution_unit_0_n_17_3),.ZN(eu_mdb_out[10]));
	AOI22_X1_LVT execution_unit_0i_13_21 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[9]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[9]),.ZN(execution_unit_0_n_13_12));
	INV_X1_LVT execution_unit_0i_13_22 (.A(execution_unit_0_n_13_12),.ZN(execution_unit_0_n_28));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b9___05F05d (.D(execution_unit_0_n_28),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(execution_unit_0_mdb_out_nxt[9]),.QN());
	AOI22_X1_LVT execution_unit_0i_13_5 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[1]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[1]),.ZN(execution_unit_0_n_13_4));
	INV_X1_LVT execution_unit_0i_13_6 (.A(execution_unit_0_n_13_4),.ZN(execution_unit_0_n_20));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b1___05F05d (.D(execution_unit_0_n_20),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(eu_mdb_out[1]),.QN());
	AOI22_X1_LVT execution_unit_0i_17_3 (.A1(execution_unit_0_n_17_0),.A2(execution_unit_0_mdb_out_nxt[9]),.B1(inst_bw),.B2(eu_mdb_out[1]),.ZN(execution_unit_0_n_17_2));
	INV_X1_LVT execution_unit_0i_17_4 (.A(execution_unit_0_n_17_2),.ZN(eu_mdb_out[9]));
	AOI22_X1_LVT execution_unit_0i_13_19 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[8]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[8]),.ZN(execution_unit_0_n_13_11));
	INV_X1_LVT execution_unit_0i_13_20 (.A(execution_unit_0_n_13_11),.ZN(execution_unit_0_n_27));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b8___05F05d (.D(execution_unit_0_n_27),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(execution_unit_0_mdb_out_nxt[8]),.QN());
	AOI22_X1_LVT execution_unit_0i_13_3 (.A1(execution_unit_0_n_13_2),.A2(execution_unit_0_alu_out[0]),.B1(execution_unit_0_n_13_1),.B2(pc_nxt[0]),.ZN(execution_unit_0_n_13_3));
	INV_X1_LVT execution_unit_0i_13_4 (.A(execution_unit_0_n_13_3),.ZN(execution_unit_0_n_19));
	DFFR_X1_LVT execution_unit_0mdb_out_nxt_reg___05F05b0___05F05d (.D(execution_unit_0_n_19),.RN(execution_unit_0_n_18),.CK(execution_unit_0_n_17),.Q(eu_mdb_out[0]),.QN());
	AOI22_X1_LVT execution_unit_0i_17_1 (.A1(execution_unit_0_n_17_0),.A2(execution_unit_0_mdb_out_nxt[8]),.B1(eu_mdb_out[0]),.B2(inst_bw),.ZN(execution_unit_0_n_17_1));
	INV_X1_LVT execution_unit_0i_17_2 (.A(execution_unit_0_n_17_1),.ZN(eu_mdb_out[8]));
	NAND3_X1_LVT clock_module_0i_7_0 (.A1(per_addr[3]),.A2(per_addr[5]),.A3(per_en),.ZN(clock_module_0_n_7_0));
	NOR4_X1_LVT clock_module_0i_7_1 (.A1(clock_module_0_n_7_0),.A2(per_addr[11]),.A3(per_addr[12]),.A4(per_addr[13]),.ZN(clock_module_0_n_7_1));
	NOR4_X1_LVT clock_module_0i_7_2 (.A1(per_addr[7]),.A2(per_addr[8]),.A3(per_addr[9]),.A4(per_addr[10]),.ZN(clock_module_0_n_7_2));
	NAND2_X1_LVT clock_module_0i_7_3 (.A1(clock_module_0_n_7_1),.A2(clock_module_0_n_7_2),.ZN(clock_module_0_n_7_3));
	NOR3_X1_LVT clock_module_0i_7_4 (.A1(clock_module_0_n_7_3),.A2(per_addr[4]),.A3(per_addr[6]),.ZN(clock_module_0_reg_sel));
	AND2_X1_LVT clock_module_0i_16_0 (.A1(per_we[1]),.A2(clock_module_0_reg_sel),.ZN(clock_module_0_reg_hi_write));
	NAND2_X1_LVT clock_module_0i_11_0 (.A1(per_addr[0]),.A2(per_addr[1]),.ZN(clock_module_0_n_11_0));
	NOR2_X1_LVT clock_module_0i_11_1 (.A1(clock_module_0_n_11_0),.A2(per_addr[2]),.ZN(clock_module_0_n_5));
	AND2_X1_LVT clock_module_0i_17_0 (.A1(clock_module_0_reg_hi_write),.A2(clock_module_0_n_5),.ZN(clock_module_0_bcsctl1_wr));
	INV_X1_LVT clock_module_0i_40_0 (.A(reset_n),.ZN(clock_module_0_por_a));
	INV_X1_LVT clock_module_0sync_cell_mclk_wkupi_0_0 (.A(puc_rst),.ZN(clock_module_0_sync_cell_mclk_wkup_n_0));
	DFFR_X1_LVT clock_module_0sync_cell_mclk_wkupdata_sync_reg___05F05b0___05F05d (.D(mclk_wkup),.RN(clock_module_0_sync_cell_mclk_wkup_n_0),.CK(dco_clk),.Q(clock_module_0_sync_cell_mclk_wkup_n_1),.QN());
	DFFR_X1_LVT clock_module_0sync_cell_mclk_wkupdata_sync_reg___05F05b1___05F05d (.D(clock_module_0_sync_cell_mclk_wkup_n_1),.RN(clock_module_0_sync_cell_mclk_wkup_n_0),.CK(dco_clk),.Q(clock_module_0_mclk_wkup_s),.QN());
	NOR2_X1_LVT clock_module_0i_37_0 (.A1(mclk_enable),.A2(clock_module_0_mclk_wkup_s),.ZN(clock_module_0_n_37_0));
	NAND2_X1_LVT clock_module_0i_37_1 (.A1(dbg_en),.A2(cpu_en),.ZN(clock_module_0_n_37_1));
	NAND2_X1_LVT clock_module_0i_37_2 (.A1(clock_module_0_n_37_0),.A2(clock_module_0_n_37_1),.ZN(clock_module_0_mclk_active));
	AND2_X1_LVT clock_module_0i_13_0 (.A1(per_we[0]),.A2(clock_module_0_reg_sel),.ZN(clock_module_0_reg_lo_write));
	INV_X1_LVT clock_module_0i_10_0 (.A(per_addr[2]),.ZN(clock_module_0_n_10_0));
	NOR3_X1_LVT clock_module_0i_10_1 (.A1(clock_module_0_n_10_0),.A2(per_addr[0]),.A3(per_addr[1]),.ZN(clock_module_0_n_4));
	AND2_X1_LVT clock_module_0i_14_0 (.A1(clock_module_0_reg_lo_write),.A2(clock_module_0_n_4),.ZN(clock_module_0_bcsctl2_wr));
	CLKGATETST_X1_LVT clock_module_0clk_gate_bcsctl2_reg (.CK(mclk),.E(clock_module_0_bcsctl2_wr),.SE(1'b0),.GCK(clock_module_0_n_8));
	DFFR_X1_LVT clock_module_0bcsctl2_reg___05F05b5___05F05d (.D(per_din[5]),.RN(clock_module_0_n_10),.CK(clock_module_0_n_8),.Q(clock_module_0_bcsctl2[5]),.QN());
	INV_X1_LVT clock_module_0i_36_2 (.A(clock_module_0_bcsctl2[5]),.ZN(clock_module_0_n_36_2));
	DFFR_X1_LVT clock_module_0bcsctl2_reg___05F05b4___05F05d (.D(per_din[4]),.RN(clock_module_0_n_10),.CK(clock_module_0_n_8),.Q(clock_module_0_bcsctl2[4]),.QN());
	OR2_X1_LVT clock_module_0i_36_3 (.A1(clock_module_0_n_36_2),.A2(clock_module_0_bcsctl2[4]),.ZN(clock_module_0_n_36_3));
	INV_X1_LVT clock_module_0i_31_0 (.A(clock_module_0_mclk_div[0]),.ZN(clock_module_0_n_19));
	OR2_X1_LVT clock_module_0i_32_0 (.A1(clock_module_0_bcsctl2[4]),.A2(clock_module_0_bcsctl2[5]),.ZN(clock_module_0_n_22));
	CLKGATETST_X1_LVT clock_module_0clk_gate_mclk_div_reg (.CK(dco_clk),.E(clock_module_0_n_22),.SE(1'b0),.GCK(clock_module_0_n_18));
	DFFR_X1_LVT clock_module_0mclk_div_reg___05F05b0___05F05d (.D(clock_module_0_n_19),.RN(clock_module_0_n_10),.CK(clock_module_0_n_18),.Q(clock_module_0_mclk_div[0]),.QN());
	HA_X1_LVT clock_module_0i_31_1 (.A(clock_module_0_mclk_div[1]),.B(clock_module_0_mclk_div[0]),.CO(clock_module_0_n_31_0),.S(clock_module_0_n_20));
	DFFR_X1_LVT clock_module_0mclk_div_reg___05F05b1___05F05d (.D(clock_module_0_n_20),.RN(clock_module_0_n_10),.CK(clock_module_0_n_18),.Q(clock_module_0_mclk_div[1]),.QN());
	XNOR2_X1_LVT clock_module_0i_31_2 (.A(clock_module_0_mclk_div[2]),.B(clock_module_0_n_31_0),.ZN(clock_module_0_n_31_1));
	INV_X1_LVT clock_module_0i_31_3 (.A(clock_module_0_n_31_1),.ZN(clock_module_0_n_21));
	DFFR_X1_LVT clock_module_0mclk_div_reg___05F05b2___05F05d (.D(clock_module_0_n_21),.RN(clock_module_0_n_10),.CK(clock_module_0_n_18),.Q(clock_module_0_mclk_div[2]),.QN());
	AND3_X1_LVT clock_module_0i_34_0 (.A1(clock_module_0_mclk_div[0]),.A2(clock_module_0_mclk_div[1]),.A3(clock_module_0_mclk_div[2]),.ZN(clock_module_0_n_23));
	INV_X1_LVT clock_module_0i_36_4 (.A(clock_module_0_n_36_3),.ZN(clock_module_0_n_36_4));
	AND2_X1_LVT clock_module_0i_35_0 (.A1(clock_module_0_mclk_div[0]),.A2(clock_module_0_mclk_div[1]),.ZN(clock_module_0_n_24));
	AOI22_X1_LVT clock_module_0i_36_5 (.A1(clock_module_0_n_36_3),.A2(clock_module_0_n_23),.B1(clock_module_0_n_36_4),.B2(clock_module_0_n_24),.ZN(clock_module_0_n_36_5));
	INV_X1_LVT clock_module_0i_36_6 (.A(clock_module_0_n_36_5),.ZN(clock_module_0_n_36_6));
	NAND2_X1_LVT clock_module_0i_36_7 (.A1(clock_module_0_n_36_2),.A2(clock_module_0_bcsctl2[4]),.ZN(clock_module_0_n_36_7));
	INV_X1_LVT clock_module_0i_36_8 (.A(clock_module_0_n_36_7),.ZN(clock_module_0_n_36_8));
	AOI22_X1_LVT clock_module_0i_36_9 (.A1(clock_module_0_n_36_6),.A2(clock_module_0_n_36_7),.B1(clock_module_0_n_36_8),.B2(clock_module_0_mclk_div[0]),.ZN(clock_module_0_n_36_9));
	NOR2_X1_LVT clock_module_0i_36_0 (.A1(clock_module_0_bcsctl2[4]),.A2(clock_module_0_bcsctl2[5]),.ZN(clock_module_0_n_36_0));
	INV_X1_LVT clock_module_0i_36_1 (.A(clock_module_0_n_36_0),.ZN(clock_module_0_n_36_1));
	NAND2_X1_LVT clock_module_0i_36_10 (.A1(clock_module_0_n_36_9),.A2(clock_module_0_n_36_1),.ZN(clock_module_0_mclk_div_sel));
	AND2_X1_LVT clock_module_0i_38_0 (.A1(clock_module_0_mclk_active),.A2(clock_module_0_mclk_div_sel),.ZN(clock_module_0_mclk_div_en));
	OR2_X1_LVT clock_module_0clock_gate_mclki_0_0 (.A1(clock_module_0_mclk_div_en),.A2(scan_enable),.ZN(clock_module_0_clock_gate_mclk_enable_in));
	INV_X1_LVT clock_module_0clock_gate_mclki_1_0 (.A(dco_clk),.ZN(clock_module_0_clock_gate_mclk_n_0));
	DLH_X1_LVT clock_module_0clock_gate_mclkenable_latch_reg (.D(clock_module_0_clock_gate_mclk_enable_in),.G(clock_module_0_clock_gate_mclk_n_0),.Q(clock_module_0_clock_gate_mclk_enable_latch));
	AND2_X1_LVT clock_module_0clock_gate_mclki_3_0 (.A1(dco_clk),.A2(clock_module_0_clock_gate_mclk_enable_latch),.ZN(cpu_mclk));
	INV_X1_LVT clock_module_0i_41_0 (.A(dbg_en),.ZN(clock_module_0_dbg_rst_nxt));
	INV_X1_LVT clock_module_0sync_reset_pori_0_0 (.A(clock_module_0_por_a),.ZN(clock_module_0_sync_reset_por_n_0));
	DFFS_X1_LVT clock_module_0sync_reset_pordata_sync_reg___05F05b0___05F05d (.D(1'b0),.SN(clock_module_0_sync_reset_por_n_0),.CK(dco_clk),.Q(clock_module_0_sync_reset_por_n_1),.QN());
	DFFS_X1_LVT clock_module_0sync_reset_pordata_sync_reg___05F05b1___05F05d (.D(clock_module_0_sync_reset_por_n_1),.SN(clock_module_0_sync_reset_por_n_0),.CK(dco_clk),.Q(clock_module_0_por_noscan),.QN());
	INV_X1_LVT clock_module_0scan_mux_pori_0_0 (.A(scan_mode),.ZN(clock_module_0_scan_mux_por_n_0_0));
	AOI22_X1_LVT clock_module_0scan_mux_pori_0_1 (.A1(clock_module_0_scan_mux_por_n_0_0),.A2(clock_module_0_por_noscan),.B1(clock_module_0_por_a),.B2(scan_mode),.ZN(clock_module_0_scan_mux_por_n_0_1));
	INV_X1_LVT clock_module_0scan_mux_pori_0_2 (.A(clock_module_0_scan_mux_por_n_0_1),.ZN(por));
	INV_X1_LVT clock_module_0i_3_0 (.A(por),.ZN(clock_module_0_n_1));
	DFFS_X1_LVT clock_module_0dbg_rst_noscan_reg (.D(clock_module_0_dbg_rst_nxt),.SN(clock_module_0_n_1),.CK(cpu_mclk),.Q(clock_module_0_dbg_rst_noscan),.QN());
	AND3_X1_LVT clock_module_0i_46_0 (.A1(dbg_en),.A2(puc_pnd_set),.A3(clock_module_0_dbg_rst_noscan),.ZN(clock_module_0_n_46_0));
	NOR2_X1_LVT clock_module_0i_46_1 (.A1(clock_module_0_n_46_0),.A2(dbg_cpu_reset),.ZN(clock_module_0_n_28));
	OR2_X1_LVT clock_module_0i_59_0 (.A1(por),.A2(wdt_reset),.ZN(clock_module_0_puc_a));
	INV_X1_LVT clock_module_0scan_mux_puc_rst_ai_0_0 (.A(scan_mode),.ZN(clock_module_0_scan_mux_puc_rst_a_n_0_0));
	AOI22_X1_LVT clock_module_0scan_mux_puc_rst_ai_0_1 (.A1(clock_module_0_scan_mux_puc_rst_a_n_0_0),.A2(clock_module_0_puc_a),.B1(clock_module_0_por_a),.B2(scan_mode),.ZN(clock_module_0_scan_mux_puc_rst_a_n_0_1));
	INV_X1_LVT clock_module_0scan_mux_puc_rst_ai_0_2 (.A(clock_module_0_scan_mux_puc_rst_a_n_0_1),.ZN(clock_module_0_puc_a_scan));
	INV_X1_LVT clock_module_0sync_cell_puci_0_0 (.A(clock_module_0_puc_a_scan),.ZN(clock_module_0_sync_cell_puc_n_0));
	DFFR_X1_LVT clock_module_0sync_cell_pucdata_sync_reg___05F05b0___05F05d (.D(clock_module_0_n_28),.RN(clock_module_0_sync_cell_puc_n_0),.CK(cpu_mclk),.Q(clock_module_0_sync_cell_puc_n_1),.QN());
	DFFR_X1_LVT clock_module_0sync_cell_pucdata_sync_reg___05F05b1___05F05d (.D(clock_module_0_sync_cell_puc_n_1),.RN(clock_module_0_sync_cell_puc_n_0),.CK(cpu_mclk),.Q(clock_module_0_puc_noscan_n),.QN());
	INV_X1_LVT clock_module_0i_21_0 (.A(clock_module_0_puc_noscan_n),.ZN(puc_pnd_set));
	INV_X1_LVT clock_module_0scan_mux_puc_rsti_0_0 (.A(scan_mode),.ZN(clock_module_0_scan_mux_puc_rst_n_0_0));
	AOI22_X1_LVT clock_module_0scan_mux_puc_rsti_0_1 (.A1(clock_module_0_scan_mux_puc_rst_n_0_0),.A2(puc_pnd_set),.B1(clock_module_0_por_a),.B2(scan_mode),.ZN(clock_module_0_scan_mux_puc_rst_n_0_1));
	INV_X1_LVT clock_module_0scan_mux_puc_rsti_0_2 (.A(clock_module_0_scan_mux_puc_rst_n_0_1),.ZN(puc_rst));
	INV_X1_LVT clock_module_0i_18_0 (.A(puc_rst),.ZN(clock_module_0_n_10));
	DFFR_X1_LVT clock_module_0bcsctl1_reg___05F05b0___05F05d (.D(per_din[8]),.RN(clock_module_0_n_10),.CK(clock_module_0_n_9),.Q(clock_module_0_bcsctl1[0]),.QN());
	AND2_X1_LVT clock_module_0and_cpuoff_mclk_dma_eni_0_0 (.A1(clock_module_0_bcsctl1[0]),.A2(mclk_dma_enable),.ZN(clock_module_0_cpuoff_and_mclk_dma_enable));
	AND2_X1_LVT clock_module_0and_cpuoff_mclk_dma_wkupi_0_0 (.A1(clock_module_0_bcsctl1[0]),.A2(mclk_dma_wkup),.ZN(clock_module_0_cpuoff_and_mclk_dma_wkup));
	INV_X1_LVT clock_module_0sync_cell_mclk_dma_wkupi_0_0 (.A(puc_rst),.ZN(clock_module_0_sync_cell_mclk_dma_wkup_n_0));
	DFFR_X1_LVT clock_module_0sync_cell_mclk_dma_wkupdata_sync_reg___05F05b0___05F05d (.D(clock_module_0_cpuoff_and_mclk_dma_wkup),.RN(clock_module_0_sync_cell_mclk_dma_wkup_n_0),.CK(dco_clk),.Q(clock_module_0_sync_cell_mclk_dma_wkup_n_1),.QN());
	DFFR_X1_LVT clock_module_0sync_cell_mclk_dma_wkupdata_sync_reg___05F05b1___05F05d (.D(clock_module_0_sync_cell_mclk_dma_wkup_n_1),.RN(clock_module_0_sync_cell_mclk_dma_wkup_n_0),.CK(dco_clk),.Q(clock_module_0_cpuoff_and_mclk_dma_wkup_s),.QN());
	OR3_X1_LVT clock_module_0i_39_0 (.A1(clock_module_0_cpuoff_and_mclk_dma_enable),.A2(clock_module_0_mclk_active),.A3(clock_module_0_cpuoff_and_mclk_dma_wkup_s),.ZN(clock_module_0_n_39_0));
	AND2_X1_LVT clock_module_0i_39_1 (.A1(clock_module_0_n_39_0),.A2(clock_module_0_mclk_div_sel),.ZN(clock_module_0_mclk_dma_div_en));
	OR2_X1_LVT clock_module_0clock_gate_dma_mclki_0_0 (.A1(clock_module_0_mclk_dma_div_en),.A2(scan_enable),.ZN(clock_module_0_clock_gate_dma_mclk_enable_in));
	INV_X1_LVT clock_module_0clock_gate_dma_mclki_1_0 (.A(dco_clk),.ZN(clock_module_0_clock_gate_dma_mclk_n_0));
	DLH_X1_LVT clock_module_0clock_gate_dma_mclkenable_latch_reg (.D(clock_module_0_clock_gate_dma_mclk_enable_in),.G(clock_module_0_clock_gate_dma_mclk_n_0),.Q(clock_module_0_clock_gate_dma_mclk_enable_latch));
	AND2_X1_LVT clock_module_0clock_gate_dma_mclki_3_0 (.A1(dco_clk),.A2(clock_module_0_clock_gate_dma_mclk_enable_latch),.ZN(mclk));
	CLKGATETST_X1_LVT clock_module_0clk_gate_bcsctl1_reg (.CK(mclk),.E(clock_module_0_bcsctl1_wr),.SE(1'b0),.GCK(clock_module_0_n_9));
	DFFR_X1_LVT clock_module_0bcsctl1_reg___05F05b5___05F05d (.D(per_din[13]),.RN(clock_module_0_n_10),.CK(clock_module_0_n_9),.Q(clock_module_0_bcsctl1[5]),.QN());
	INV_X1_LVT clock_module_0i_28_2 (.A(clock_module_0_bcsctl1[5]),.ZN(clock_module_0_n_28_2));
	DFFR_X1_LVT clock_module_0bcsctl1_reg___05F05b4___05F05d (.D(per_din[12]),.RN(clock_module_0_n_10),.CK(clock_module_0_n_9),.Q(clock_module_0_bcsctl1[4]),.QN());
	OR2_X1_LVT clock_module_0i_28_3 (.A1(clock_module_0_n_28_2),.A2(clock_module_0_bcsctl1[4]),.ZN(clock_module_0_n_28_3));
	INV_X1_LVT clock_module_0i_23_0 (.A(clock_module_0_aclk_div[0]),.ZN(clock_module_0_n_12));
	OR2_X1_LVT clock_module_0i_24_0 (.A1(clock_module_0_bcsctl1[4]),.A2(clock_module_0_bcsctl1[5]),.ZN(clock_module_0_n_15));
	CLKGATETST_X1_LVT clock_module_0clk_gate_aclk_div_reg (.CK(dco_clk),.E(clock_module_0_n_15),.SE(1'b0),.GCK(clock_module_0_n_11));
	DFFR_X1_LVT clock_module_0aclk_div_reg___05F05b0___05F05d (.D(clock_module_0_n_12),.RN(clock_module_0_n_10),.CK(clock_module_0_n_11),.Q(clock_module_0_aclk_div[0]),.QN());
	HA_X1_LVT clock_module_0i_23_1 (.A(clock_module_0_aclk_div[1]),.B(clock_module_0_aclk_div[0]),.CO(clock_module_0_n_23_0),.S(clock_module_0_n_13));
	DFFR_X1_LVT clock_module_0aclk_div_reg___05F05b1___05F05d (.D(clock_module_0_n_13),.RN(clock_module_0_n_10),.CK(clock_module_0_n_11),.Q(clock_module_0_aclk_div[1]),.QN());
	XNOR2_X1_LVT clock_module_0i_23_2 (.A(clock_module_0_aclk_div[2]),.B(clock_module_0_n_23_0),.ZN(clock_module_0_n_23_1));
	INV_X1_LVT clock_module_0i_23_3 (.A(clock_module_0_n_23_1),.ZN(clock_module_0_n_14));
	DFFR_X1_LVT clock_module_0aclk_div_reg___05F05b2___05F05d (.D(clock_module_0_n_14),.RN(clock_module_0_n_10),.CK(clock_module_0_n_11),.Q(clock_module_0_aclk_div[2]),.QN());
	AND3_X1_LVT clock_module_0i_26_0 (.A1(clock_module_0_aclk_div[0]),.A2(clock_module_0_aclk_div[1]),.A3(clock_module_0_aclk_div[2]),.ZN(clock_module_0_n_16));
	INV_X1_LVT clock_module_0i_28_4 (.A(clock_module_0_n_28_3),.ZN(clock_module_0_n_28_4));
	AND2_X1_LVT clock_module_0i_27_0 (.A1(clock_module_0_aclk_div[0]),.A2(clock_module_0_aclk_div[1]),.ZN(clock_module_0_n_17));
	AOI22_X1_LVT clock_module_0i_28_5 (.A1(clock_module_0_n_28_3),.A2(clock_module_0_n_16),.B1(clock_module_0_n_28_4),.B2(clock_module_0_n_17),.ZN(clock_module_0_n_28_5));
	INV_X1_LVT clock_module_0i_28_6 (.A(clock_module_0_n_28_5),.ZN(clock_module_0_n_28_6));
	NAND2_X1_LVT clock_module_0i_28_7 (.A1(clock_module_0_n_28_2),.A2(clock_module_0_bcsctl1[4]),.ZN(clock_module_0_n_28_7));
	INV_X1_LVT clock_module_0i_28_8 (.A(clock_module_0_n_28_7),.ZN(clock_module_0_n_28_8));
	AOI22_X1_LVT clock_module_0i_28_9 (.A1(clock_module_0_n_28_6),.A2(clock_module_0_n_28_7),.B1(clock_module_0_n_28_8),.B2(clock_module_0_aclk_div[0]),.ZN(clock_module_0_n_28_9));
	NOR2_X1_LVT clock_module_0i_28_0 (.A1(clock_module_0_bcsctl1[4]),.A2(clock_module_0_bcsctl1[5]),.ZN(clock_module_0_n_28_0));
	INV_X1_LVT clock_module_0i_28_1 (.A(clock_module_0_n_28_0),.ZN(clock_module_0_n_28_1));
	NAND2_X1_LVT clock_module_0i_28_10 (.A1(clock_module_0_n_28_9),.A2(clock_module_0_n_28_1),.ZN(clock_module_0_aclk_div_sel));
	NAND2_X1_LVT clock_module_0i_29_0 (.A1(cpu_en),.A2(clock_module_0_aclk_div_sel),.ZN(clock_module_0_n_29_0));
	NOR2_X1_LVT clock_module_0i_29_1 (.A1(clock_module_0_n_29_0),.A2(oscoff),.ZN(clock_module_0_aclk_div_en));
	OR2_X1_LVT clock_module_0clock_gate_aclki_0_0 (.A1(clock_module_0_aclk_div_en),.A2(scan_enable),.ZN(clock_module_0_clock_gate_aclk_enable_in));
	INV_X1_LVT clock_module_0clock_gate_aclki_1_0 (.A(dco_clk),.ZN(clock_module_0_clock_gate_aclk_n_0));
	DLH_X1_LVT clock_module_0clock_gate_aclkenable_latch_reg (.D(clock_module_0_clock_gate_aclk_enable_in),.G(clock_module_0_clock_gate_aclk_n_0),.Q(clock_module_0_clock_gate_aclk_enable_latch));
	AND2_X1_LVT clock_module_0clock_gate_aclki_3_0 (.A1(dco_clk),.A2(clock_module_0_clock_gate_aclk_enable_latch),.ZN(aclk));
	OR2_X1_LVT clock_module_0clock_gate_dbg_clki_0_0 (.A1(dbg_en),.A2(scan_enable),.ZN(clock_module_0_clock_gate_dbg_clk_enable_in));
	INV_X1_LVT clock_module_0clock_gate_dbg_clki_1_0 (.A(cpu_mclk),.ZN(clock_module_0_clock_gate_dbg_clk_n_0));
	DLH_X1_LVT clock_module_0clock_gate_dbg_clkenable_latch_reg (.D(clock_module_0_clock_gate_dbg_clk_enable_in),.G(clock_module_0_clock_gate_dbg_clk_n_0),.Q(clock_module_0_clock_gate_dbg_clk_enable_latch));
	AND2_X1_LVT clock_module_0clock_gate_dbg_clki_3_0 (.A1(cpu_mclk),.A2(clock_module_0_clock_gate_dbg_clk_enable_latch),.ZN(dbg_clk));
	INV_X1_LVT clock_module_0scan_mux_dbg_rsti_0_0 (.A(scan_mode),.ZN(clock_module_0_scan_mux_dbg_rst_n_0_0));
	AOI22_X1_LVT clock_module_0scan_mux_dbg_rsti_0_1 (.A1(clock_module_0_scan_mux_dbg_rst_n_0_0),.A2(clock_module_0_dbg_rst_noscan),.B1(clock_module_0_por_a),.B2(scan_mode),.ZN(clock_module_0_scan_mux_dbg_rst_n_0_1));
	INV_X1_LVT clock_module_0scan_mux_dbg_rsti_0_2 (.A(clock_module_0_scan_mux_dbg_rst_n_0_1),.ZN(dbg_rst));
	DFFR_X1_LVT clock_module_0bcsctl2_reg___05F05b7___05F05d (.D(1'b0),.RN(clock_module_0_n_10),.CK(clock_module_0_n_8),.Q(clock_module_0_bcsctl2[7]),.QN());
	INV_X1_LVT clock_module_0i_58_0 (.A(clock_module_0_bcsctl2[7]),.ZN(clock_module_0_n_39));
	AND2_X1_LVT clock_module_0and_dco_mclk_wkupi_0_0 (.A1(mclk_wkup),.A2(clock_module_0_n_39),.ZN(clock_module_0_dco_mclk_wkup));
	INV_X1_LVT clock_module_0i_57_0 (.A(dco_enable),.ZN(clock_module_0_n_38));
	AND2_X1_LVT clock_module_0and_cpuoff_mclk_eni_0_0 (.A1(cpuoff),.A2(mclk_enable),.ZN(clock_module_0_cpuoff_and_mclk_enable));
	AND2_X1_LVT clock_module_0and_dco_dis1i_0_0 (.A1(clock_module_0_n_39),.A2(clock_module_0_cpuoff_and_mclk_enable),.ZN(clock_module_0_cpu_enabled_with_dco));
	DFFR_X1_LVT clock_module_0bcsctl1_reg___05F05b2___05F05d (.D(per_din[10]),.RN(clock_module_0_n_10),.CK(clock_module_0_n_9),.Q(clock_module_0_bcsctl1[2]),.QN());
	AND2_X1_LVT clock_module_0and_scg0_mclk_dma_eni_0_0 (.A1(clock_module_0_bcsctl1[2]),.A2(mclk_dma_enable),.ZN(clock_module_0_scg0_and_mclk_dma_enable));
	NOR2_X1_LVT clock_module_0i_60_0 (.A1(clock_module_0_cpu_enabled_with_dco),.A2(clock_module_0_scg0_and_mclk_dma_enable),.ZN(clock_module_0_n_40));
	AND2_X1_LVT clock_module_0and_dco_dis2i_0_0 (.A1(clock_module_0_dbg_rst_nxt),.A2(clock_module_0_n_40),.ZN(clock_module_0_dco_not_enabled_by_dbg));
	AND2_X1_LVT clock_module_0and_dco_dis3i_0_0 (.A1(scg0),.A2(clock_module_0_dco_not_enabled_by_dbg),.ZN(clock_module_0_dco_disable_by_scg0));
	INV_X1_LVT clock_module_0i_42_0 (.A(clock_module_0_dco_disable_by_scg0),.ZN(clock_module_0_n_25));
	INV_X1_LVT clock_module_0i_55_0 (.A(cpu_en),.ZN(clock_module_0_n_36));
	INV_X1_LVT clock_module_0i_56_0 (.A(mclk_enable),.ZN(clock_module_0_n_37));
	AND2_X1_LVT clock_module_0and_dco_dis4i_0_0 (.A1(clock_module_0_n_36),.A2(clock_module_0_n_37),.ZN(clock_module_0_dco_disable_by_cpu_en));
	INV_X1_LVT clock_module_0i_43_0 (.A(clock_module_0_dco_disable_by_cpu_en),.ZN(clock_module_0_n_26));
	AND2_X1_LVT clock_module_0and_dco_dis5i_0_0 (.A1(clock_module_0_n_25),.A2(clock_module_0_n_26),.ZN(clock_module_0_dco_enable_nxt));
	AND2_X1_LVT clock_module_0and_dco_en_wkupi_0_0 (.A1(clock_module_0_n_38),.A2(clock_module_0_dco_enable_nxt),.ZN(clock_module_0_dco_en_wkup));
	AND2_X1_LVT clock_module_0and_scg0_mclk_dma_wkupi_0_0 (.A1(clock_module_0_bcsctl1[2]),.A2(mclk_dma_wkup),.ZN(clock_module_0_scg0_and_mclk_dma_wkup));
	OR3_X1_LVT clock_module_0i_44_0 (.A1(clock_module_0_dco_mclk_wkup),.A2(clock_module_0_dco_en_wkup),.A3(clock_module_0_scg0_and_mclk_dma_wkup),.ZN(clock_module_0_dco_wkup_set));
	INV_X1_LVT clock_module_0scan_mux_dco_wkup_observei_0_0 (.A(scan_mode),.ZN(clock_module_0_scan_mux_dco_wkup_observe_n_0_0));
	AOI22_X1_LVT clock_module_0scan_mux_dco_wkup_observei_0_1 (.A1(clock_module_0_scan_mux_dco_wkup_observe_n_0_0),.A2(1'b0),.B1(clock_module_0_dco_wkup_set),.B2(scan_mode),.ZN(clock_module_0_scan_mux_dco_wkup_observe_n_0_1));
	INV_X1_LVT clock_module_0scan_mux_dco_wkup_observei_0_2 (.A(clock_module_0_scan_mux_dco_wkup_observe_n_0_1),.ZN(clock_module_0_dco_wkup_set_scan_observe));
	INV_X1_LVT clock_module_0i_1_0 (.A(clock_module_0_dco_wkup_set_scan_observe),.ZN(clock_module_0_n_1_0));
	NAND2_X1_LVT clock_module_0i_1_1 (.A1(clock_module_0_n_1_0),.A2(clock_module_0_dco_enable_nxt),.ZN(clock_module_0_n_0));
	DFFS_X1_LVT clock_module_0dco_disable_reg (.D(clock_module_0_n_0),.SN(clock_module_0_n_1),.CK(dco_clk),.Q(clock_module_0_dco_disable),.QN());
	INV_X1_LVT clock_module_0i_5_0 (.A(clock_module_0_dco_disable),.ZN(clock_module_0_n_2));
	INV_X1_LVT clock_module_0i_0_0 (.A(dco_clk),.ZN(clock_module_0_nodiv_mclk_n));
	DFFR_X1_LVT clock_module_0dco_enable_reg (.D(clock_module_0_n_2),.RN(clock_module_0_n_1),.CK(clock_module_0_nodiv_mclk_n),.Q(dco_enable),.QN());
	OR2_X1_LVT clock_module_0i_61_0 (.A1(clock_module_0_dco_wkup_set),.A2(por),.ZN(clock_module_0_n_41));
	INV_X1_LVT clock_module_0scan_mux_dco_wkupi_0_0 (.A(scan_mode),.ZN(clock_module_0_scan_mux_dco_wkup_n_0_0));
	AOI22_X1_LVT clock_module_0scan_mux_dco_wkupi_0_1 (.A1(clock_module_0_scan_mux_dco_wkup_n_0_0),.A2(clock_module_0_n_41),.B1(clock_module_0_por_a),.B2(scan_mode),.ZN(clock_module_0_scan_mux_dco_wkup_n_0_1));
	INV_X1_LVT clock_module_0scan_mux_dco_wkupi_0_2 (.A(clock_module_0_scan_mux_dco_wkup_n_0_1),.ZN(clock_module_0_dco_wkup_set_scan));
	INV_X1_LVT clock_module_0sync_cell_dco_wkupi_0_0 (.A(clock_module_0_dco_wkup_set_scan),.ZN(clock_module_0_sync_cell_dco_wkup_n_0));
	DFFR_X1_LVT clock_module_0sync_cell_dco_wkupdata_sync_reg___05F05b0___05F05d (.D(1'b1),.RN(clock_module_0_sync_cell_dco_wkup_n_0),.CK(clock_module_0_nodiv_mclk_n),.Q(clock_module_0_sync_cell_dco_wkup_n_1),.QN());
	DFFR_X1_LVT clock_module_0sync_cell_dco_wkupdata_sync_reg___05F05b1___05F05d (.D(clock_module_0_sync_cell_dco_wkup_n_1),.RN(clock_module_0_sync_cell_dco_wkup_n_0),.CK(clock_module_0_nodiv_mclk_n),.Q(clock_module_0_dco_wkup_n),.QN());
	INV_X1_LVT clock_module_0i_45_0 (.A(clock_module_0_dco_wkup_n),.ZN(clock_module_0_n_27));
	AND2_X1_LVT clock_module_0and_dco_wkupi_0_0 (.A1(clock_module_0_n_27),.A2(cpu_en),.ZN(dco_wkup));
	NOR2_X1_LVT clock_module_0i_8_0 (.A1(per_we[0]),.A2(per_we[1]),.ZN(clock_module_0_n_3));
	AND2_X1_LVT clock_module_0i_9_0 (.A1(clock_module_0_n_3),.A2(clock_module_0_reg_sel),.ZN(clock_module_0_reg_read));
	AND2_X1_LVT clock_module_0i_12_0 (.A1(clock_module_0_reg_read),.A2(clock_module_0_n_5),.ZN(clock_module_0_n_6));
	DFFR_X1_LVT clock_module_0bcsctl1_reg___05F05b7___05F05d (.D(1'b0),.RN(clock_module_0_n_10),.CK(clock_module_0_n_9),.Q(clock_module_0_bcsctl1[7]),.QN());
	AND2_X1_LVT clock_module_0i_20_15 (.A1(clock_module_0_n_6),.A2(clock_module_0_bcsctl1[7]),.ZN(per_dout_clk[15]));
	DFFR_X1_LVT clock_module_0bcsctl1_reg___05F05b6___05F05d (.D(1'b0),.RN(clock_module_0_n_10),.CK(clock_module_0_n_9),.Q(clock_module_0_bcsctl1[6]),.QN());
	AND2_X1_LVT clock_module_0i_20_14 (.A1(clock_module_0_n_6),.A2(clock_module_0_bcsctl1[6]),.ZN(per_dout_clk[14]));
	AND2_X1_LVT clock_module_0i_20_13 (.A1(clock_module_0_n_6),.A2(clock_module_0_bcsctl1[5]),.ZN(per_dout_clk[13]));
	AND2_X1_LVT clock_module_0i_20_12 (.A1(clock_module_0_n_6),.A2(clock_module_0_bcsctl1[4]),.ZN(per_dout_clk[12]));
	DFFR_X1_LVT clock_module_0bcsctl1_reg___05F05b3___05F05d (.D(per_din[11]),.RN(clock_module_0_n_10),.CK(clock_module_0_n_9),.Q(clock_module_0_bcsctl1[3]),.QN());
	AND2_X1_LVT clock_module_0i_20_11 (.A1(clock_module_0_n_6),.A2(clock_module_0_bcsctl1[3]),.ZN(per_dout_clk[11]));
	AND2_X1_LVT clock_module_0i_20_10 (.A1(clock_module_0_n_6),.A2(clock_module_0_bcsctl1[2]),.ZN(per_dout_clk[10]));
	DFFR_X1_LVT clock_module_0bcsctl1_reg___05F05b1___05F05d (.D(1'b0),.RN(clock_module_0_n_10),.CK(clock_module_0_n_9),.Q(clock_module_0_bcsctl1[1]),.QN());
	AND2_X1_LVT clock_module_0i_20_9 (.A1(clock_module_0_n_6),.A2(clock_module_0_bcsctl1[1]),.ZN(per_dout_clk[9]));
	AND2_X1_LVT clock_module_0i_20_8 (.A1(clock_module_0_bcsctl1[0]),.A2(clock_module_0_n_6),.ZN(per_dout_clk[8]));
	AND2_X1_LVT clock_module_0i_12_1 (.A1(clock_module_0_reg_read),.A2(clock_module_0_n_4),.ZN(clock_module_0_n_7));
	AND2_X1_LVT clock_module_0i_20_7 (.A1(clock_module_0_n_7),.A2(clock_module_0_bcsctl2[7]),.ZN(per_dout_clk[7]));
	DFFR_X1_LVT clock_module_0bcsctl2_reg___05F05b6___05F05d (.D(1'b0),.RN(clock_module_0_n_10),.CK(clock_module_0_n_8),.Q(clock_module_0_bcsctl2[6]),.QN());
	AND2_X1_LVT clock_module_0i_20_6 (.A1(clock_module_0_n_7),.A2(clock_module_0_bcsctl2[6]),.ZN(per_dout_clk[6]));
	AND2_X1_LVT clock_module_0i_20_5 (.A1(clock_module_0_n_7),.A2(clock_module_0_bcsctl2[5]),.ZN(per_dout_clk[5]));
	AND2_X1_LVT clock_module_0i_20_4 (.A1(clock_module_0_n_7),.A2(clock_module_0_bcsctl2[4]),.ZN(per_dout_clk[4]));
	DFFR_X1_LVT clock_module_0bcsctl2_reg___05F05b3___05F05d (.D(1'b0),.RN(clock_module_0_n_10),.CK(clock_module_0_n_8),.Q(clock_module_0_bcsctl2[3]),.QN());
	AND2_X1_LVT clock_module_0i_20_3 (.A1(clock_module_0_n_7),.A2(clock_module_0_bcsctl2[3]),.ZN(per_dout_clk[3]));
	DFFR_X1_LVT clock_module_0bcsctl2_reg___05F05b2___05F05d (.D(per_din[2]),.RN(clock_module_0_n_10),.CK(clock_module_0_n_8),.Q(clock_module_0_bcsctl2[2]),.QN());
	AND2_X1_LVT clock_module_0i_20_2 (.A1(clock_module_0_n_7),.A2(clock_module_0_bcsctl2[2]),.ZN(per_dout_clk[2]));
	DFFR_X1_LVT clock_module_0bcsctl2_reg___05F05b1___05F05d (.D(per_din[1]),.RN(clock_module_0_n_10),.CK(clock_module_0_n_8),.Q(clock_module_0_bcsctl2[1]),.QN());
	AND2_X1_LVT clock_module_0i_20_1 (.A1(clock_module_0_n_7),.A2(clock_module_0_bcsctl2[1]),.ZN(per_dout_clk[1]));
	DFFR_X1_LVT clock_module_0bcsctl2_reg___05F05b0___05F05d (.D(1'b0),.RN(clock_module_0_n_10),.CK(clock_module_0_n_8),.Q(clock_module_0_bcsctl2[0]),.QN());
	AND2_X1_LVT clock_module_0i_20_0 (.A1(clock_module_0_bcsctl2[0]),.A2(clock_module_0_n_7),.ZN(per_dout_clk[0]));
	INV_X1_LVT clock_module_0i_54_0 (.A(scg1),.ZN(clock_module_0_n_54_0));
	AND2_X1_LVT clock_module_0and_scg1_mclk_dma_wkupi_0_0 (.A1(clock_module_0_bcsctl1[3]),.A2(mclk_dma_wkup),.ZN(clock_module_0_scg1_and_mclk_dma_wkup));
	INV_X1_LVT clock_module_0sync_cell_smclk_dma_wkupi_0_0 (.A(puc_rst),.ZN(clock_module_0_sync_cell_smclk_dma_wkup_n_0));
	DFFR_X1_LVT clock_module_0sync_cell_smclk_dma_wkupdata_sync_reg___05F05b0___05F05d (.D(clock_module_0_scg1_and_mclk_dma_wkup),.RN(clock_module_0_sync_cell_smclk_dma_wkup_n_0),.CK(dco_clk),.Q(clock_module_0_sync_cell_smclk_dma_wkup_n_1),.QN());
	DFFR_X1_LVT clock_module_0sync_cell_smclk_dma_wkupdata_sync_reg___05F05b1___05F05d (.D(clock_module_0_sync_cell_smclk_dma_wkup_n_1),.RN(clock_module_0_sync_cell_smclk_dma_wkup_n_0),.CK(dco_clk),.Q(clock_module_0_scg1_and_mclk_dma_wkup_s),.QN());
	AND2_X1_LVT clock_module_0and_scg1_mclk_dma_eni_0_0 (.A1(clock_module_0_bcsctl1[3]),.A2(mclk_dma_enable),.ZN(clock_module_0_scg1_and_mclk_dma_enable));
	NOR3_X1_LVT clock_module_0i_54_1 (.A1(clock_module_0_n_54_0),.A2(clock_module_0_scg1_and_mclk_dma_wkup_s),.A3(clock_module_0_scg1_and_mclk_dma_enable),.ZN(clock_module_0_n_54_1));
	INV_X1_LVT clock_module_0i_53_2 (.A(clock_module_0_bcsctl2[2]),.ZN(clock_module_0_n_53_2));
	OR2_X1_LVT clock_module_0i_53_3 (.A1(clock_module_0_n_53_2),.A2(clock_module_0_bcsctl2[1]),.ZN(clock_module_0_n_53_3));
	INV_X1_LVT clock_module_0i_48_0 (.A(clock_module_0_smclk_div[0]),.ZN(clock_module_0_n_30));
	OR2_X1_LVT clock_module_0i_49_0 (.A1(clock_module_0_bcsctl2[1]),.A2(clock_module_0_bcsctl2[2]),.ZN(clock_module_0_n_33));
	CLKGATETST_X1_LVT clock_module_0clk_gate_smclk_div_reg (.CK(dco_clk),.E(clock_module_0_n_33),.SE(1'b0),.GCK(clock_module_0_n_29));
	DFFR_X1_LVT clock_module_0smclk_div_reg___05F05b0___05F05d (.D(clock_module_0_n_30),.RN(clock_module_0_n_10),.CK(clock_module_0_n_29),.Q(clock_module_0_smclk_div[0]),.QN());
	HA_X1_LVT clock_module_0i_48_1 (.A(clock_module_0_smclk_div[1]),.B(clock_module_0_smclk_div[0]),.CO(clock_module_0_n_48_0),.S(clock_module_0_n_31));
	DFFR_X1_LVT clock_module_0smclk_div_reg___05F05b1___05F05d (.D(clock_module_0_n_31),.RN(clock_module_0_n_10),.CK(clock_module_0_n_29),.Q(clock_module_0_smclk_div[1]),.QN());
	XNOR2_X1_LVT clock_module_0i_48_2 (.A(clock_module_0_smclk_div[2]),.B(clock_module_0_n_48_0),.ZN(clock_module_0_n_48_1));
	INV_X1_LVT clock_module_0i_48_3 (.A(clock_module_0_n_48_1),.ZN(clock_module_0_n_32));
	DFFR_X1_LVT clock_module_0smclk_div_reg___05F05b2___05F05d (.D(clock_module_0_n_32),.RN(clock_module_0_n_10),.CK(clock_module_0_n_29),.Q(clock_module_0_smclk_div[2]),.QN());
	AND3_X1_LVT clock_module_0i_51_0 (.A1(clock_module_0_smclk_div[0]),.A2(clock_module_0_smclk_div[1]),.A3(clock_module_0_smclk_div[2]),.ZN(clock_module_0_n_34));
	INV_X1_LVT clock_module_0i_53_4 (.A(clock_module_0_n_53_3),.ZN(clock_module_0_n_53_4));
	AND2_X1_LVT clock_module_0i_52_0 (.A1(clock_module_0_smclk_div[0]),.A2(clock_module_0_smclk_div[1]),.ZN(clock_module_0_n_35));
	AOI22_X1_LVT clock_module_0i_53_5 (.A1(clock_module_0_n_53_3),.A2(clock_module_0_n_34),.B1(clock_module_0_n_53_4),.B2(clock_module_0_n_35),.ZN(clock_module_0_n_53_5));
	INV_X1_LVT clock_module_0i_53_6 (.A(clock_module_0_n_53_5),.ZN(clock_module_0_n_53_6));
	NAND2_X1_LVT clock_module_0i_53_7 (.A1(clock_module_0_n_53_2),.A2(clock_module_0_bcsctl2[1]),.ZN(clock_module_0_n_53_7));
	INV_X1_LVT clock_module_0i_53_8 (.A(clock_module_0_n_53_7),.ZN(clock_module_0_n_53_8));
	AOI22_X1_LVT clock_module_0i_53_9 (.A1(clock_module_0_n_53_6),.A2(clock_module_0_n_53_7),.B1(clock_module_0_n_53_8),.B2(clock_module_0_smclk_div[0]),.ZN(clock_module_0_n_53_9));
	NOR2_X1_LVT clock_module_0i_53_0 (.A1(clock_module_0_bcsctl2[1]),.A2(clock_module_0_bcsctl2[2]),.ZN(clock_module_0_n_53_0));
	INV_X1_LVT clock_module_0i_53_1 (.A(clock_module_0_n_53_0),.ZN(clock_module_0_n_53_1));
	NAND2_X1_LVT clock_module_0i_53_10 (.A1(clock_module_0_n_53_9),.A2(clock_module_0_n_53_1),.ZN(clock_module_0_smclk_div_sel));
	NAND2_X1_LVT clock_module_0i_54_2 (.A1(cpu_en),.A2(clock_module_0_smclk_div_sel),.ZN(clock_module_0_n_54_2));
	NOR2_X1_LVT clock_module_0i_54_3 (.A1(clock_module_0_n_54_1),.A2(clock_module_0_n_54_2),.ZN(clock_module_0_smclk_div_en));
	OR2_X1_LVT clock_module_0clock_gate_smclki_0_0 (.A1(clock_module_0_smclk_div_en),.A2(scan_enable),.ZN(clock_module_0_clock_gate_smclk_enable_in));
	INV_X1_LVT clock_module_0clock_gate_smclki_1_0 (.A(dco_clk),.ZN(clock_module_0_clock_gate_smclk_n_0));
	DLH_X1_LVT clock_module_0clock_gate_smclkenable_latch_reg (.D(clock_module_0_clock_gate_smclk_enable_in),.G(clock_module_0_clock_gate_smclk_n_0),.Q(clock_module_0_clock_gate_smclk_enable_latch));
	AND2_X1_LVT clock_module_0clock_gate_smclki_3_0 (.A1(dco_clk),.A2(clock_module_0_clock_gate_smclk_enable_latch),.ZN(smclk));
endmodule