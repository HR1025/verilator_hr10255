module DFFR_X1_LVT(Q,QN,CK,D,RN);
	 output Q;
	 output QN;
	 input CK;
	 input D;
	 input RN;


endmodule

module AOI22_X1_LVT(ZN,A1,A2,B1,B2);
	 output ZN;
	 input A1;
	 input A2;
	 input B1;
	 input B2;


endmodule

module OAI22_X1_LVT(ZN,A1,A2,B1,B2);
	 output ZN;
	 input A1;
	 input A2;
	 input B1;
	 input B2;


endmodule

module NOR4_X1_LVT(ZN,A1,A2,A3,A4);
	 output ZN;
	 input A1;
	 input A2;
	 input A3;
	 input A4;


endmodule

module NOR3_X1_LVT(ZN,A1,A2,A3);
	 output ZN;
	 input A1;
	 input A2;
	 input A3;


endmodule

module XNOR2_X1_LVT(ZN,A,B);
	 output ZN;
	 input A;
	 input B;


endmodule

module OR2_X1_LVT(ZN,A1,A2);
	 output ZN;
	 input A1;
	 input A2;


endmodule

module OAI211_X1_LVT(ZN,A,B,C1,C2);
	 output ZN;
	 input A;
	 input B;
	 input C1;
	 input C2;


endmodule

module NAND4_X1_LVT(ZN,A1,A2,A3,A4);
	 output ZN;
	 input A1;
	 input A2;
	 input A3;
	 input A4;


endmodule

module HA_X1_LVT(CO,S,A,B);
	 output CO;
	 output S;
	 input A;
	 input B;


endmodule

module NAND3_X1_LVT(ZN,A1,A2,A3);
	 output ZN;
	 input A1;
	 input A2;
	 input A3;


endmodule

module FA_X1_LVT(CO,S,A,B,CI);
	 output CO;
	 output S;
	 input A;
	 input B;
	 input CI;


endmodule

module DLH_X1_LVT(Q,D,G);
	 output Q;
	 input D;
	 input G;


endmodule

module CLKGATETST_X1_LVT(GCK,CK,E,SE);
	 output GCK;
	 input CK;
	 input E;
	 input SE;


endmodule

module AOI222_X1_LVT(ZN,A1,A2,B1,B2,C1,C2);
	 output ZN;
	 input A1;
	 input A2;
	 input B1;
	 input B2;
	 input C1;
	 input C2;


endmodule

module AOI21_X1_LVT(ZN,A,B1,B2);
	 output ZN;
	 input A;
	 input B1;
	 input B2;


endmodule

module AOI211_X1_LVT(ZN,A,B,C1,C2);
	 output ZN;
	 input A;
	 input B;
	 input C1;
	 input C2;


endmodule

module omsp_sync_cell(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_scan_mux(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module OAI33_X1_LVT(ZN,A1,A2,A3,B1,B2,B3);
	 output ZN;
	 input A1;
	 input A2;
	 input A3;
	 input B1;
	 input B2;
	 input B3;


endmodule

module OAI21_X1_LVT(ZN,A,B1,B2);
	 output ZN;
	 input A;
	 input B1;
	 input B2;


endmodule

module omsp_clock_gate(gclk,clk,enable,scan_enable);
	 output gclk;
	 input clk;
	 input enable;
	 input scan_enable;

	 wire enable_in;
	 wire enable_latch;
	 wire n_0;

endmodule

module omsp_and_gate__2_57(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_and_gate__2_53(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_sync_cell__2_23(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module INV_X1_LVT(ZN,A);
	 output ZN;
	 input A;


endmodule

module AND3_X1_LVT(ZN,A1,A2,A3);
	 output ZN;
	 input A1;
	 input A2;
	 input A3;


endmodule

module omsp_scan_mux__2_67(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module DFFS_X1_LVT(Q,QN,CK,D,SN);
	 output Q;
	 output QN;
	 input CK;
	 input D;
	 input SN;


endmodule

module omsp_and_gate__1_5(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_and_gate__1_1(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_scan_mux__2_69(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module omsp_sync_cell__2_17(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_sync_cell__2_27(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_and_gate__0_1424(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module AOI221_X1_LVT(ZN,A,B1,B2,C1,C2);
	 output ZN;
	 input A;
	 input B1;
	 input B2;
	 input C1;
	 input C2;


endmodule

module omsp_and_gate__2_41(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_and_gate(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_execution_unit(cpuoff,dbg_reg_din,gie,mab,mb_en,mb_wr,mdb_out,oscoff,pc_sw,pc_sw_wr,scg0,scg1,dbg_halt_st,dbg_mem_dout,dbg_reg_wr,e_state,exec_done,inst_ad,inst_as,inst_alu,inst_bw,inst_dest,inst_dext,inst_irq_rst,inst_jmp,inst_mov,inst_sext,inst_so,inst_src,inst_type,mclk,mdb_in,pc,pc_nxt,puc_rst,scan_enable);
	 output cpuoff;
	 output [15:0]dbg_reg_din;
	 output gie;
	 output [15:0]mab;
	 output mb_en;
	 output [1:0]mb_wr;
	 output [15:0]mdb_out;
	 output oscoff;
	 output [15:0]pc_sw;
	 output pc_sw_wr;
	 output scg0;
	 output scg1;
	 input dbg_halt_st;
	 input [15:0]dbg_mem_dout;
	 input dbg_reg_wr;
	 input [3:0]e_state;
	 input exec_done;
	 input [7:0]inst_ad;
	 input [7:0]inst_as;
	 input [11:0]inst_alu;
	 input inst_bw;
	 input [15:0]inst_dest;
	 input [15:0]inst_dext;
	 input inst_irq_rst;
	 input [7:0]inst_jmp;
	 input inst_mov;
	 input [15:0]inst_sext;
	 input [7:0]inst_so;
	 input [15:0]inst_src;
	 input [2:0]inst_type;
	 input mclk;
	 input [15:0]mdb_in;
	 input [15:0]pc;
	 input [15:0]pc_nxt;
	 input puc_rst;
	 input scan_enable;

	 wire [3:0]alu_stat_wr;
	 wire [3:0]alu_stat;
	 wire [15:0]alu_out;
	 wire [3:0]status;
	 wire [15:0]reg_src;
	 wire n_0_0;
	 wire n_0_1;
	 wire n_0_2;
	 wire n_0_3;
	 wire reg_sr_clr;
	 wire n_4_0;
	 wire n_4_1;
	 wire mb_wr_det;
	 wire n_7_0;
	 wire n_7_1;
	 wire n_7_2;
	 wire n_7_3;
	 wire n_7_4;
	 wire n_8_0;
	 wire n_8_1;
	 wire n_8_2;
	 wire n_8_3;
	 wire mab_lsb;
	 wire [15:0]mdb_out_nxt;
	 wire n_13_0;
	 wire n_13_1;
	 wire n_13_2;
	 wire n_13_3;
	 wire n_13_4;
	 wire n_13_5;
	 wire n_13_6;
	 wire n_13_7;
	 wire n_13_8;
	 wire n_13_9;
	 wire n_13_10;
	 wire n_13_11;
	 wire n_13_12;
	 wire n_13_13;
	 wire n_13_14;
	 wire n_13_15;
	 wire n_13_16;
	 wire n_13_17;
	 wire n_13_18;
	 wire n_14_0;
	 wire n_14_1;
	 wire n_15_0;
	 wire n_15_1;
	 wire n_15_2;
	 wire n_15_3;
	 wire n_17_0;
	 wire n_17_1;
	 wire n_17_2;
	 wire n_17_3;
	 wire n_17_4;
	 wire n_17_5;
	 wire n_17_6;
	 wire n_17_7;
	 wire n_17_8;
	 wire n_21_0;
	 wire n_21_1;
	 wire n_21_2;
	 wire n_21_3;
	 wire n_21_4;
	 wire reg_dest_wr;
	 wire n_23_0;
	 wire reg_pc_call;
	 wire n_30_0;
	 wire n_30_1;
	 wire n_30_2;
	 wire reg_sp_wr;
	 wire reg_sr_wr;
	 wire n_32_0;
	 wire reg_incr;
	 wire n_34_0;
	 wire n_34_1;
	 wire n_34_2;
	 wire n_34_3;
	 wire n_34_4;
	 wire n_34_5;
	 wire n_34_6;
	 wire n_34_7;
	 wire n_34_8;
	 wire n_34_9;
	 wire n_34_10;
	 wire n_34_11;
	 wire n_34_12;
	 wire n_34_13;
	 wire n_34_14;
	 wire n_34_15;
	 wire n_34_16;
	 wire n_34_17;
	 wire n_39_0;
	 wire n_39_1;
	 wire n_39_2;
	 wire n_39_3;
	 wire n_39_4;
	 wire n_39_5;
	 wire n_39_6;
	 wire n_39_7;
	 wire n_39_8;
	 wire n_40_0;
	 wire n_40_1;
	 wire n_40_2;
	 wire n_40_3;
	 wire n_40_4;
	 wire n_40_5;
	 wire n_40_6;
	 wire n_41_0;
	 wire n_41_1;
	 wire n_41_2;
	 wire n_41_3;
	 wire n_41_4;
	 wire n_41_5;
	 wire n_41_6;
	 wire n_41_7;
	 wire n_41_8;
	 wire n_41_9;
	 wire n_41_10;
	 wire n_41_11;
	 wire n_41_12;
	 wire n_41_13;
	 wire n_41_14;
	 wire n_41_15;
	 wire n_41_16;
	 wire n_41_17;
	 wire n_41_18;
	 wire n_41_19;
	 wire n_41_20;
	 wire n_41_21;
	 wire n_41_22;
	 wire n_41_23;
	 wire n_41_24;
	 wire n_41_25;
	 wire n_41_26;
	 wire n_41_27;
	 wire n_41_28;
	 wire n_41_29;
	 wire n_41_30;
	 wire n_41_31;
	 wire n_41_32;
	 wire n_41_33;
	 wire n_41_34;
	 wire n_41_35;
	 wire n_41_36;
	 wire n_41_37;
	 wire n_41_38;
	 wire n_41_39;
	 wire n_41_40;
	 wire n_41_41;
	 wire n_41_42;
	 wire n_41_43;
	 wire n_41_44;
	 wire n_41_45;
	 wire n_41_46;
	 wire n_41_47;
	 wire n_41_48;
	 wire n_41_49;
	 wire n_41_50;
	 wire n_41_51;
	 wire n_41_52;
	 wire n_41_53;
	 wire n_41_54;
	 wire n_41_55;
	 wire n_41_56;
	 wire n_41_57;
	 wire n_41_58;
	 wire n_41_59;
	 wire n_41_60;
	 wire n_41_61;
	 wire n_41_62;
	 wire n_41_63;
	 wire n_41_64;
	 wire n_41_65;
	 wire n_41_66;
	 wire n_41_67;
	 wire n_41_68;
	 wire n_41_69;
	 wire n_41_70;
	 wire n_41_71;
	 wire n_41_72;
	 wire n_41_73;
	 wire n_41_74;
	 wire n_41_75;
	 wire n_41_76;
	 wire n_41_77;
	 wire n_41_78;
	 wire n_41_79;
	 wire mdb_in_buf_en;
	 wire [15:0]mdb_in_buf;
	 wire mdb_in_buf_valid;
	 wire n_44_0;
	 wire n_44_1;
	 wire n_45_0;
	 wire n_45_1;
	 wire n_45_2;
	 wire n_48_0;
	 wire n_48_1;
	 wire n_48_2;
	 wire n_48_3;
	 wire n_48_4;
	 wire n_48_5;
	 wire n_48_6;
	 wire n_48_7;
	 wire n_48_8;
	 wire n_48_9;
	 wire n_49_0;
	 wire n_49_1;
	 wire n_49_2;
	 wire n_49_3;
	 wire n_49_4;
	 wire n_49_5;
	 wire n_49_6;
	 wire n_49_7;
	 wire n_49_8;
	 wire n_49_9;
	 wire n_50_0;
	 wire n_50_1;
	 wire n_50_2;
	 wire n_50_3;
	 wire n_50_4;
	 wire n_50_5;
	 wire n_50_6;
	 wire n_50_7;
	 wire n_50_8;
	 wire n_50_9;
	 wire n_50_10;
	 wire n_50_11;
	 wire n_50_12;
	 wire n_50_13;
	 wire n_50_14;
	 wire n_50_15;
	 wire n_50_16;
	 wire n_50_17;
	 wire n_50_18;
	 wire n_50_19;
	 wire n_50_20;
	 wire n_50_21;
	 wire n_50_22;
	 wire n_50_23;
	 wire n_50_24;
	 wire n_50_25;
	 wire n_50_26;
	 wire n_50_27;
	 wire n_50_28;
	 wire n_50_29;
	 wire n_50_30;
	 wire n_50_31;
	 wire n_50_32;
	 wire n_50_33;
	 wire n_50_34;
	 wire n_50_35;
	 wire n_50_36;
	 wire n_50_37;
	 wire n_50_38;
	 wire n_50_39;
	 wire n_50_40;
	 wire n_50_41;
	 wire n_50_42;
	 wire n_50_43;
	 wire n_50_44;
	 wire n_50_45;
	 wire n_50_46;
	 wire n_50_47;
	 wire n_50_48;
	 wire n_50_49;
	 wire n_50_50;
	 wire n_50_51;
	 wire n_50_52;
	 wire n_50_53;
	 wire n_50_54;
	 wire n_50_55;
	 wire n_50_56;
	 wire n_50_57;
	 wire n_50_58;
	 wire n_50_59;
	 wire n_50_60;
	 wire n_50_61;
	 wire n_50_62;
	 wire n_50_63;
	 wire n_50_64;
	 wire n_50_65;
	 wire n_50_66;
	 wire n_50_67;
	 wire n_50_68;
	 wire n_50_69;
	 wire n_50_70;
	 wire n_50_71;
	 wire n_50_72;
	 wire n_50_73;
	 wire n_50_74;
	 wire n_50_75;
	 wire n_50_76;
	 wire n_50_77;
	 wire n_50_78;
	 wire n_50_79;
	 wire n_50_80;
	 wire n_50_81;
	 wire n_50_82;
	 wire n_50_83;
	 wire n_50_84;
	 wire n_50_85;
	 wire n_50_86;
	 wire n_50_87;
	 wire n_50_88;
	 wire n_50_89;
	 wire n_50_90;
	 wire n_50_91;
	 wire n_50_92;
	 wire n_50_93;
	 wire n_50_94;
	 wire n_50_95;
	 wire n_0;
	 wire n_69;
	 wire n_1;
	 wire n_2;
	 wire n_73;
	 wire n_74;
	 wire n_3;
	 wire n_40;
	 wire n_10;
	 wire n_67;
	 wire n_68;
	 wire n_72;
	 wire n_75;
	 wire n_47;
	 wire n_13;
	 wire n_11;
	 wire n_6;
	 wire n_5;
	 wire n_12;
	 wire n_4;
	 wire n_9;
	 wire n_16;
	 wire n_18;
	 wire n_49;
	 wire n_48;
	 wire n_65;
	 wire n_37;
	 wire n_38;
	 wire n_71;
	 wire n_76;
	 wire n_41;
	 wire n_42;
	 wire n_43;
	 wire n_8;
	 wire n_44;
	 wire n_46;
	 wire n_66;
	 wire n_7;
	 wire n_45;
	 wire n_70;
	 wire n_77;
	 wire n_93;
	 wire n_64;
	 wire n_92;
	 wire n_63;
	 wire n_91;
	 wire n_62;
	 wire n_90;
	 wire n_61;
	 wire n_89;
	 wire n_60;
	 wire n_88;
	 wire n_59;
	 wire n_87;
	 wire n_58;
	 wire n_86;
	 wire n_57;
	 wire n_85;
	 wire n_56;
	 wire n_84;
	 wire n_55;
	 wire n_83;
	 wire n_54;
	 wire n_82;
	 wire n_53;
	 wire n_81;
	 wire n_52;
	 wire n_80;
	 wire n_51;
	 wire n_79;
	 wire n_50;
	 wire n_78;
	 wire n_102;
	 wire n_98;
	 wire n_103;
	 wire n_96;
	 wire n_97;
	 wire n_95;
	 wire n_101;
	 wire n_105;
	 wire n_94;
	 wire n_106;
	 wire n_39;
	 wire n_100;
	 wire n_107;
	 wire n_99;
	 wire n_108;
	 wire n_104;
	 wire n_124;
	 wire n_123;
	 wire n_122;
	 wire n_121;
	 wire n_120;
	 wire n_119;
	 wire n_118;
	 wire n_117;
	 wire n_116;
	 wire n_115;
	 wire n_114;
	 wire n_113;
	 wire n_112;
	 wire n_111;
	 wire n_110;
	 wire n_109;
	 wire n_15;
	 wire n_14;
	 wire n_34;
	 wire n_35;
	 wire n_36;
	 wire n_17;
	 wire n_26;
	 wire n_33;
	 wire n_25;
	 wire n_32;
	 wire n_24;
	 wire n_31;
	 wire n_23;
	 wire n_30;
	 wire n_22;
	 wire n_29;
	 wire n_21;
	 wire n_28;
	 wire n_20;
	 wire n_27;
	 wire n_19;

endmodule

module AND2_X1_LVT(ZN,A1,A2);
	 output ZN;
	 input A1;
	 input A2;


endmodule

module omsp_sync_cell__0_1430(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_scan_mux__2_71(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module omsp_scan_mux__2_63(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module omsp_scan_mux__2_59(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module omsp_clock_module(aclk,aclk_en,cpu_en_s,cpu_mclk,dma_mclk,dbg_clk,dbg_en_s,dbg_rst,dco_enable,dco_wkup,lfxt_enable,lfxt_wkup,per_dout,por,puc_pnd_set,puc_rst,smclk,smclk_en,cpu_en,cpuoff,dbg_cpu_reset,dbg_en,dco_clk,lfxt_clk,mclk_dma_enable,mclk_dma_wkup,mclk_enable,mclk_wkup,oscoff,per_addr,per_din,per_en,per_we,reset_n,scan_enable,scan_mode,scg0,scg1,wdt_reset);
	 output aclk;
	 output aclk_en;
	 output cpu_en_s;
	 output cpu_mclk;
	 output dma_mclk;
	 output dbg_clk;
	 output dbg_en_s;
	 output dbg_rst;
	 output dco_enable;
	 output dco_wkup;
	 output lfxt_enable;
	 output lfxt_wkup;
	 output [15:0]per_dout;
	 output por;
	 output puc_pnd_set;
	 output puc_rst;
	 output smclk;
	 output smclk_en;
	 input cpu_en;
	 input cpuoff;
	 input dbg_cpu_reset;
	 input dbg_en;
	 input dco_clk;
	 input lfxt_clk;
	 input mclk_dma_enable;
	 input mclk_dma_wkup;
	 input mclk_enable;
	 input mclk_wkup;
	 input oscoff;
	 input [13:0]per_addr;
	 input [15:0]per_din;
	 input per_en;
	 input [1:0]per_we;
	 input reset_n;
	 input scan_enable;
	 input scan_mode;
	 input scg0;
	 input scg1;
	 input wdt_reset;

	 wire cpuoff_and_mclk_dma_wkup;
	 wire cpuoff_and_mclk_dma_wkup_s;
	 wire mclk_wkup_s;
	 wire cpuoff_and_mclk_dma_enable;
	 wire por_noscan;
	 wire puc_a_scan;
	 wire puc_noscan_n;
	 wire scg0_and_mclk_dma_enable;
	 wire cpuoff_and_mclk_enable;
	 wire cpu_enabled_with_dco;
	 wire dco_not_enabled_by_dbg;
	 wire dco_disable_by_scg0;
	 wire dco_disable_by_cpu_en;
	 wire dco_enable_nxt;
	 wire scg0_and_mclk_dma_wkup;
	 wire dco_en_wkup;
	 wire dco_mclk_wkup;
	 wire dco_wkup_set_scan_observe;
	 wire dco_wkup_set_scan;
	 wire dco_wkup_n;
	 wire scg1_and_mclk_dma_enable;
	 wire scg1_and_mclk_dma_wkup;
	 wire scg1_and_mclk_dma_wkup_s;
	 wire nodiv_mclk_n;
	 wire dco_disable;
	 wire n_1_0;
	 wire n_7_0;
	 wire n_7_1;
	 wire n_7_2;
	 wire n_7_3;
	 wire reg_sel;
	 wire reg_read;
	 wire n_10_0;
	 wire n_11_0;
	 wire reg_lo_write;
	 wire bcsctl2_wr;
	 wire [7:0]bcsctl2;
	 wire reg_hi_write;
	 wire bcsctl1_wr;
	 wire [7:0]bcsctl1;
	 wire [2:0]aclk_div;
	 wire n_23_0;
	 wire n_23_1;
	 wire n_28_0;
	 wire n_28_1;
	 wire n_28_2;
	 wire n_28_3;
	 wire n_28_4;
	 wire n_28_5;
	 wire n_28_6;
	 wire n_28_7;
	 wire n_28_8;
	 wire n_28_9;
	 wire aclk_div_sel;
	 wire n_29_0;
	 wire aclk_div_en;
	 wire [2:0]mclk_div;
	 wire n_31_0;
	 wire n_31_1;
	 wire n_36_0;
	 wire n_36_1;
	 wire n_36_2;
	 wire n_36_3;
	 wire n_36_4;
	 wire n_36_5;
	 wire n_36_6;
	 wire n_36_7;
	 wire n_36_8;
	 wire n_36_9;
	 wire mclk_div_sel;
	 wire n_37_0;
	 wire n_37_1;
	 wire mclk_active;
	 wire mclk_div_en;
	 wire n_39_0;
	 wire mclk_dma_div_en;
	 wire por_a;
	 wire dbg_rst_nxt;
	 wire dbg_rst_noscan;
	 wire dco_wkup_set;
	 wire n_46_0;
	 wire [2:0]smclk_div;
	 wire n_48_0;
	 wire n_48_1;
	 wire n_53_0;
	 wire n_53_1;
	 wire n_53_2;
	 wire n_53_3;
	 wire n_53_4;
	 wire n_53_5;
	 wire n_53_6;
	 wire n_53_7;
	 wire n_53_8;
	 wire n_53_9;
	 wire smclk_div_sel;
	 wire n_54_0;
	 wire n_54_1;
	 wire n_54_2;
	 wire smclk_div_en;
	 wire puc_a;
	 wire n_5;
	 wire n_4;
	 wire n_8;
	 wire n_10;
	 wire n_19;
	 wire n_22;
	 wire n_18;
	 wire n_20;
	 wire n_21;
	 wire n_23;
	 wire n_24;
	 wire n_1;
	 wire n_28;
	 wire n_9;
	 wire n_12;
	 wire n_15;
	 wire n_11;
	 wire n_13;
	 wire n_14;
	 wire n_16;
	 wire n_17;
	 wire n_39;
	 wire n_38;
	 wire n_40;
	 wire n_25;
	 wire n_36;
	 wire n_37;
	 wire n_26;
	 wire n_0;
	 wire n_2;
	 wire n_41;
	 wire n_27;
	 wire n_3;
	 wire n_6;
	 wire n_7;
	 wire n_30;
	 wire n_33;
	 wire n_29;
	 wire n_31;
	 wire n_32;
	 wire n_34;
	 wire n_35;

endmodule

module NAND2_X1_LVT(ZN,A1,A2);
	 output ZN;
	 input A1;
	 input A2;


endmodule

module omsp_watchdog(per_dout,wdt_irq,wdt_reset,wdt_wkup,wdtifg,wdtnmies,aclk,aclk_en,dbg_freeze,mclk,per_addr,per_din,per_en,per_we,por,puc_rst,scan_enable,scan_mode,smclk,smclk_en,wdtie,wdtifg_irq_clr,wdtifg_sw_clr,wdtifg_sw_set);
	 output [15:0]per_dout;
	 output wdt_irq;
	 output wdt_reset;
	 output wdt_wkup;
	 output wdtifg;
	 output wdtnmies;
	 input aclk;
	 input aclk_en;
	 input dbg_freeze;
	 input mclk;
	 input [13:0]per_addr;
	 input [15:0]per_din;
	 input per_en;
	 input [1:0]per_we;
	 input por;
	 input puc_rst;
	 input scan_enable;
	 input scan_mode;
	 input smclk;
	 input smclk_en;
	 input wdtie;
	 input wdtifg_irq_clr;
	 input wdtifg_sw_clr;
	 input wdtifg_sw_set;

	 wire wdt_rst_noscan;
	 wire wdt_rst;
	 wire wdtcnt_incr;
	 wire wdtcnt_clr_sync;
	 wire wdt_evt_toggle_sync;
	 wire wdt_wkup_pre;
	 wire n_0_0;
	 wire n_0_1;
	 wire n_0_2;
	 wire n_0_3;
	 wire n_0_4;
	 wire reg_wr;
	 wire [7:0]wdtctl;
	 wire n_8_0;
	 wire n_8_1;
	 wire n_8_2;
	 wire wdtpw_error;
	 wire wdt_evt_toggle_sync_dly;
	 wire n_9_0;
	 wire wdtifg_set;
	 wire n_10_0;
	 wire wdtifg_clr;
	 wire n_13_0;
	 wire n_13_1;
	 wire n_17_0;
	 wire wdtcnt_clr_sync_dly;
	 wire n_19_0;
	 wire wdtcnt_clr;
	 wire [15:0]wdtcnt;
	 wire n_21_0;
	 wire n_22_0;
	 wire n_22_1;
	 wire [15:0]wdtcnt_nxt;
	 wire n_24_0;
	 wire n_24_1;
	 wire n_24_2;
	 wire n_24_3;
	 wire n_24_4;
	 wire n_24_5;
	 wire n_24_6;
	 wire n_24_7;
	 wire n_24_8;
	 wire n_24_9;
	 wire n_24_10;
	 wire n_24_11;
	 wire n_24_12;
	 wire n_24_13;
	 wire n_24_14;
	 wire [1:0]wdtisx_ss;
	 wire [1:0]wdtisx_s;
	 wire n_28_0;
	 wire n_28_1;
	 wire n_28_2;
	 wire n_28_3;
	 wire n_28_4;
	 wire n_28_5;
	 wire n_28_6;
	 wire n_28_7;
	 wire n_28_8;
	 wire wdtqn_reg;
	 wire wdtqn_edge;
	 wire wdt_evt_toggle;
	 wire wdt_wkup_en;
	 wire n_35_0;
	 wire n_35_1;
	 wire n_37_0;
	 wire wdtcnt_clr_detect;
	 wire wdtcnt_clr_toggle;
	 wire wdtifg_clr_reg;
	 wire wdtqn_edge_reg;
	 wire n_1;
	 wire n_0;
	 wire n_2;
	 wire n_3;
	 wire n_4;
	 wire n_30;
	 wire n_29;
	 wire n_35;
	 wire n_34;
	 wire n_17;
	 wire n_31;
	 wire n_33;
	 wire n_27;
	 wire n_10;
	 wire n_16;
	 wire n_15;
	 wire n_14;
	 wire n_13;
	 wire n_12;
	 wire n_11;
	 wire n_26;
	 wire n_25;
	 wire n_24;
	 wire n_23;
	 wire n_22;
	 wire n_21;
	 wire n_20;
	 wire n_19;
	 wire n_18;
	 wire n_28;
	 wire n_7;
	 wire n_5;
	 wire n_6;
	 wire n_8;
	 wire n_9;
	 wire n_32;

	assign per_dout[15] = 1'b0;
	assign per_dout[14] = per_dout[5];
	assign per_dout[13] = per_dout[5];
	assign per_dout[12] = 1'b0;
	assign per_dout[11] = per_dout[5];
	assign per_dout[9] = 1'b0;
	assign per_dout[10] = 1'b1;
	assign per_dout[8] = per_dout[5];
endmodule

module omsp_sync_cell__1_11(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_wakeup_cell__0_1428(wkup_out,scan_clk,scan_mode,scan_rst,wkup_clear,wkup_event);
	 output wkup_out;
	 input scan_clk;
	 input scan_mode;
	 input scan_rst;
	 input wkup_clear;
	 input wkup_event;

	 wire wkup_rst;
	 wire wkup_clk;
	 wire n_0;

endmodule

module omsp_scan_mux__0_1427(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module omsp_multiplier(per_dout,mclk,per_addr,per_din,per_en,per_we,puc_rst,scan_enable);
	 output [15:0]per_dout;
	 input mclk;
	 input [13:0]per_addr;
	 input [15:0]per_din;
	 input per_en;
	 input [1:0]per_we;
	 input puc_rst;
	 input scan_enable;

	 wire n_0_0;
	 wire n_0_1;
	 wire n_0_2;
	 wire n_0_3;
	 wire reg_sel;
	 wire reg_read;
	 wire n_3_0;
	 wire n_3_1;
	 wire n_3_2;
	 wire reg_rd1;
	 wire reg_rd15;
	 wire reg_write;
	 wire op2_wr;
	 wire reslo_wr;
	 wire reshi_wr;
	 wire [15:0]per_din_msk;
	 wire [15:0]op2_reg;
	 wire [1:0]cycle;
	 wire result_wr;
	 wire op1_wr;
	 wire sign_sel;
	 wire [8:0]op2_hi_xp;
	 wire n_29_0;
	 wire n_29_1;
	 wire [8:0]op2_xp;
	 wire n_29_2;
	 wire n_29_3;
	 wire n_29_4;
	 wire n_29_5;
	 wire n_29_6;
	 wire n_29_7;
	 wire n_29_8;
	 wire [15:0]op1;
	 wire [16:0]op1_xp;
	 wire n_32_0;
	 wire n_32_1;
	 wire n_32_2;
	 wire n_32_3;
	 wire n_32_4;
	 wire n_32_5;
	 wire n_32_6;
	 wire n_32_7;
	 wire n_32_8;
	 wire n_32_9;
	 wire n_32_10;
	 wire n_32_11;
	 wire n_32_12;
	 wire n_32_13;
	 wire n_32_14;
	 wire n_32_15;
	 wire n_32_16;
	 wire n_32_17;
	 wire n_32_18;
	 wire n_32_19;
	 wire n_32_20;
	 wire n_32_21;
	 wire n_32_22;
	 wire n_32_23;
	 wire n_32_24;
	 wire n_32_25;
	 wire n_32_26;
	 wire n_32_27;
	 wire n_32_28;
	 wire n_32_29;
	 wire n_32_30;
	 wire n_32_31;
	 wire n_32_32;
	 wire n_32_33;
	 wire n_32_34;
	 wire n_32_35;
	 wire n_32_36;
	 wire n_32_37;
	 wire n_32_38;
	 wire n_32_39;
	 wire n_32_40;
	 wire n_32_41;
	 wire n_32_42;
	 wire n_32_43;
	 wire n_32_44;
	 wire n_32_45;
	 wire n_32_46;
	 wire n_32_47;
	 wire n_32_48;
	 wire n_32_49;
	 wire n_32_50;
	 wire n_32_51;
	 wire n_32_52;
	 wire n_32_53;
	 wire n_32_54;
	 wire n_32_55;
	 wire n_32_56;
	 wire n_32_57;
	 wire n_32_58;
	 wire n_32_59;
	 wire n_32_60;
	 wire n_32_61;
	 wire n_32_62;
	 wire n_32_63;
	 wire n_32_64;
	 wire n_32_65;
	 wire n_32_66;
	 wire n_32_67;
	 wire n_32_68;
	 wire n_32_69;
	 wire n_32_70;
	 wire n_32_71;
	 wire n_32_72;
	 wire n_32_73;
	 wire n_32_74;
	 wire n_32_75;
	 wire n_32_76;
	 wire n_32_77;
	 wire n_32_78;
	 wire n_32_79;
	 wire n_32_80;
	 wire n_32_81;
	 wire n_32_82;
	 wire n_32_83;
	 wire n_32_84;
	 wire n_32_85;
	 wire n_32_86;
	 wire n_32_87;
	 wire n_32_88;
	 wire n_32_89;
	 wire n_32_90;
	 wire n_32_91;
	 wire n_32_92;
	 wire n_32_93;
	 wire n_32_94;
	 wire n_32_95;
	 wire n_32_96;
	 wire n_32_97;
	 wire n_32_98;
	 wire n_32_99;
	 wire n_32_100;
	 wire n_32_101;
	 wire n_32_102;
	 wire n_32_103;
	 wire n_32_104;
	 wire n_32_105;
	 wire n_32_106;
	 wire n_32_107;
	 wire n_32_108;
	 wire n_32_109;
	 wire n_32_110;
	 wire n_32_111;
	 wire n_32_112;
	 wire n_32_113;
	 wire n_32_114;
	 wire n_32_115;
	 wire n_32_116;
	 wire n_32_117;
	 wire n_32_118;
	 wire n_32_119;
	 wire n_32_120;
	 wire n_32_121;
	 wire n_32_122;
	 wire n_32_123;
	 wire n_32_124;
	 wire n_32_125;
	 wire n_32_126;
	 wire n_32_127;
	 wire n_32_128;
	 wire n_32_129;
	 wire n_32_130;
	 wire n_32_131;
	 wire n_32_132;
	 wire n_32_133;
	 wire n_32_134;
	 wire n_32_135;
	 wire n_32_136;
	 wire n_32_137;
	 wire n_32_138;
	 wire n_32_139;
	 wire n_32_140;
	 wire n_32_141;
	 wire n_32_142;
	 wire n_32_143;
	 wire n_32_144;
	 wire n_32_145;
	 wire n_32_146;
	 wire n_32_147;
	 wire n_32_148;
	 wire n_32_149;
	 wire n_32_150;
	 wire n_32_151;
	 wire n_32_152;
	 wire n_32_153;
	 wire n_32_154;
	 wire n_32_155;
	 wire n_32_156;
	 wire n_32_157;
	 wire n_32_158;
	 wire n_32_159;
	 wire n_32_160;
	 wire n_32_161;
	 wire n_32_162;
	 wire n_32_163;
	 wire n_32_164;
	 wire n_32_165;
	 wire n_32_166;
	 wire n_32_167;
	 wire n_32_168;
	 wire n_32_169;
	 wire n_32_170;
	 wire n_32_171;
	 wire n_32_172;
	 wire n_32_173;
	 wire n_32_174;
	 wire n_32_175;
	 wire n_32_176;
	 wire n_32_177;
	 wire n_32_178;
	 wire n_32_179;
	 wire n_32_180;
	 wire n_32_181;
	 wire n_32_182;
	 wire n_32_183;
	 wire n_32_184;
	 wire n_32_185;
	 wire n_32_186;
	 wire n_32_187;
	 wire n_32_188;
	 wire n_32_189;
	 wire n_32_190;
	 wire n_32_191;
	 wire n_32_192;
	 wire n_32_193;
	 wire n_32_194;
	 wire n_32_195;
	 wire n_32_196;
	 wire n_32_197;
	 wire n_32_198;
	 wire n_32_199;
	 wire n_32_200;
	 wire n_32_201;
	 wire n_32_202;
	 wire n_32_203;
	 wire n_32_204;
	 wire n_32_205;
	 wire n_32_206;
	 wire n_32_207;
	 wire n_32_208;
	 wire n_32_209;
	 wire n_32_210;
	 wire n_32_211;
	 wire n_32_212;
	 wire n_32_213;
	 wire n_32_214;
	 wire n_32_215;
	 wire n_32_216;
	 wire n_32_217;
	 wire n_32_218;
	 wire n_32_219;
	 wire n_32_220;
	 wire n_32_221;
	 wire n_32_222;
	 wire n_32_223;
	 wire n_32_224;
	 wire n_32_225;
	 wire n_32_226;
	 wire n_32_227;
	 wire n_32_228;
	 wire n_32_229;
	 wire n_32_230;
	 wire n_32_231;
	 wire n_32_232;
	 wire n_32_233;
	 wire n_32_234;
	 wire n_32_235;
	 wire n_32_236;
	 wire n_32_237;
	 wire n_32_238;
	 wire n_32_239;
	 wire n_32_240;
	 wire n_32_241;
	 wire n_32_242;
	 wire n_32_243;
	 wire n_32_244;
	 wire n_32_245;
	 wire n_32_246;
	 wire n_32_247;
	 wire n_32_248;
	 wire n_32_249;
	 wire n_32_250;
	 wire n_32_251;
	 wire n_32_252;
	 wire n_32_253;
	 wire n_32_254;
	 wire n_32_255;
	 wire n_32_256;
	 wire n_32_257;
	 wire n_32_258;
	 wire n_32_259;
	 wire n_32_260;
	 wire n_32_261;
	 wire n_32_262;
	 wire n_32_263;
	 wire n_32_264;
	 wire n_32_265;
	 wire n_32_266;
	 wire n_32_267;
	 wire n_32_268;
	 wire n_32_269;
	 wire n_32_270;
	 wire n_32_271;
	 wire n_32_272;
	 wire n_32_273;
	 wire n_32_274;
	 wire n_32_275;
	 wire n_32_276;
	 wire n_32_277;
	 wire n_32_278;
	 wire n_32_279;
	 wire n_32_280;
	 wire n_32_281;
	 wire n_32_282;
	 wire n_32_283;
	 wire n_32_284;
	 wire n_32_285;
	 wire n_32_286;
	 wire n_32_287;
	 wire n_32_288;
	 wire n_32_289;
	 wire n_32_290;
	 wire n_32_291;
	 wire n_32_292;
	 wire n_32_293;
	 wire n_32_294;
	 wire n_32_295;
	 wire n_32_296;
	 wire n_32_297;
	 wire n_32_298;
	 wire n_32_299;
	 wire n_32_300;
	 wire n_32_301;
	 wire n_32_302;
	 wire n_32_303;
	 wire n_32_304;
	 wire n_32_305;
	 wire n_32_306;
	 wire n_32_307;
	 wire n_32_308;
	 wire n_32_309;
	 wire n_32_310;
	 wire n_32_311;
	 wire n_32_312;
	 wire n_32_313;
	 wire n_32_314;
	 wire n_32_315;
	 wire n_32_316;
	 wire n_32_317;
	 wire n_32_318;
	 wire n_32_319;
	 wire n_32_320;
	 wire n_32_321;
	 wire n_32_322;
	 wire n_32_323;
	 wire n_32_324;
	 wire n_32_325;
	 wire n_32_326;
	 wire n_32_327;
	 wire n_32_328;
	 wire n_32_329;
	 wire n_32_330;
	 wire n_32_331;
	 wire n_32_332;
	 wire n_32_333;
	 wire n_32_334;
	 wire n_32_335;
	 wire n_32_336;
	 wire n_32_337;
	 wire n_32_338;
	 wire n_32_339;
	 wire n_32_340;
	 wire n_32_341;
	 wire n_32_342;
	 wire n_32_343;
	 wire n_32_344;
	 wire n_32_345;
	 wire n_32_346;
	 wire n_32_347;
	 wire n_32_348;
	 wire n_32_349;
	 wire n_32_350;
	 wire n_32_351;
	 wire n_32_352;
	 wire n_32_353;
	 wire n_32_354;
	 wire n_32_355;
	 wire n_32_356;
	 wire n_32_357;
	 wire n_32_358;
	 wire n_32_359;
	 wire n_32_360;
	 wire n_32_361;
	 wire n_32_362;
	 wire n_32_363;
	 wire n_32_364;
	 wire n_32_365;
	 wire n_32_366;
	 wire n_32_367;
	 wire n_32_368;
	 wire n_32_369;
	 wire n_32_370;
	 wire n_32_371;
	 wire n_32_372;
	 wire n_32_373;
	 wire n_32_374;
	 wire n_32_375;
	 wire n_32_376;
	 wire n_32_377;
	 wire n_32_378;
	 wire n_32_379;
	 wire n_32_380;
	 wire n_32_381;
	 wire n_32_382;
	 wire n_32_383;
	 wire n_32_384;
	 wire n_32_385;
	 wire n_32_386;
	 wire n_32_387;
	 wire n_32_388;
	 wire n_32_389;
	 wire n_32_390;
	 wire n_32_391;
	 wire n_32_392;
	 wire n_32_393;
	 wire n_32_394;
	 wire n_32_395;
	 wire n_32_396;
	 wire n_32_397;
	 wire n_32_398;
	 wire n_32_399;
	 wire n_32_400;
	 wire n_32_401;
	 wire n_32_402;
	 wire n_32_403;
	 wire n_32_404;
	 wire n_32_405;
	 wire n_32_406;
	 wire n_32_407;
	 wire n_32_408;
	 wire n_32_409;
	 wire n_32_410;
	 wire n_32_411;
	 wire n_32_412;
	 wire n_32_413;
	 wire n_32_414;
	 wire n_32_415;
	 wire n_32_416;
	 wire n_32_417;
	 wire n_32_418;
	 wire n_32_419;
	 wire n_32_420;
	 wire n_32_421;
	 wire n_32_422;
	 wire n_32_423;
	 wire n_32_424;
	 wire n_32_425;
	 wire n_32_426;
	 wire n_32_427;
	 wire n_32_428;
	 wire n_32_429;
	 wire n_32_430;
	 wire n_32_431;
	 wire n_32_432;
	 wire n_32_433;
	 wire n_32_434;
	 wire n_32_435;
	 wire n_32_436;
	 wire n_32_437;
	 wire n_32_438;
	 wire n_32_439;
	 wire n_32_440;
	 wire n_32_441;
	 wire n_32_442;
	 wire n_32_443;
	 wire n_32_444;
	 wire n_32_445;
	 wire n_32_446;
	 wire n_32_447;
	 wire n_32_448;
	 wire n_32_449;
	 wire n_32_450;
	 wire n_32_451;
	 wire n_32_452;
	 wire n_32_453;
	 wire n_32_454;
	 wire n_32_455;
	 wire n_32_456;
	 wire n_32_457;
	 wire n_32_458;
	 wire n_32_459;
	 wire n_32_460;
	 wire n_32_461;
	 wire n_32_462;
	 wire n_32_463;
	 wire n_32_464;
	 wire n_32_465;
	 wire n_32_466;
	 wire n_32_467;
	 wire n_32_468;
	 wire n_32_469;
	 wire n_32_470;
	 wire n_32_471;
	 wire n_32_472;
	 wire n_32_473;
	 wire n_32_474;
	 wire n_32_475;
	 wire n_32_476;
	 wire n_32_477;
	 wire n_32_478;
	 wire n_32_479;
	 wire n_32_480;
	 wire n_32_481;
	 wire n_32_482;
	 wire n_32_483;
	 wire n_32_484;
	 wire n_32_485;
	 wire n_32_486;
	 wire n_32_487;
	 wire n_32_488;
	 wire n_32_489;
	 wire n_32_490;
	 wire n_32_491;
	 wire n_32_492;
	 wire n_32_493;
	 wire n_32_494;
	 wire n_32_495;
	 wire n_32_496;
	 wire n_32_497;
	 wire n_32_498;
	 wire n_32_499;
	 wire n_32_500;
	 wire n_32_501;
	 wire n_32_502;
	 wire n_32_503;
	 wire n_32_504;
	 wire n_32_505;
	 wire n_32_506;
	 wire n_32_507;
	 wire n_32_508;
	 wire n_32_509;
	 wire n_32_510;
	 wire n_32_511;
	 wire n_32_512;
	 wire n_32_513;
	 wire n_32_514;
	 wire n_32_515;
	 wire n_32_516;
	 wire n_32_517;
	 wire n_32_518;
	 wire n_32_519;
	 wire n_32_520;
	 wire n_32_521;
	 wire n_32_522;
	 wire n_32_523;
	 wire n_32_524;
	 wire n_32_525;
	 wire n_32_526;
	 wire n_32_527;
	 wire n_32_528;
	 wire n_32_529;
	 wire n_32_530;
	 wire n_32_531;
	 wire n_32_532;
	 wire n_32_533;
	 wire n_32_534;
	 wire n_32_535;
	 wire n_32_536;
	 wire n_32_537;
	 wire n_32_538;
	 wire n_32_539;
	 wire n_32_540;
	 wire n_32_541;
	 wire n_32_542;
	 wire n_32_543;
	 wire n_32_544;
	 wire n_32_545;
	 wire n_32_546;
	 wire n_32_547;
	 wire n_32_548;
	 wire n_32_549;
	 wire n_32_550;
	 wire n_32_551;
	 wire n_32_552;
	 wire n_32_553;
	 wire n_32_554;
	 wire n_32_555;
	 wire n_32_556;
	 wire n_32_557;
	 wire n_32_558;
	 wire n_32_559;
	 wire n_32_560;
	 wire n_32_561;
	 wire n_32_562;
	 wire n_32_563;
	 wire n_32_564;
	 wire n_32_565;
	 wire n_32_566;
	 wire n_32_567;
	 wire n_32_568;
	 wire n_32_569;
	 wire n_32_570;
	 wire n_32_571;
	 wire n_32_572;
	 wire n_32_573;
	 wire n_32_574;
	 wire n_32_575;
	 wire n_32_576;
	 wire n_32_577;
	 wire n_32_578;
	 wire n_32_579;
	 wire n_32_580;
	 wire n_32_581;
	 wire n_32_582;
	 wire n_32_583;
	 wire n_32_584;
	 wire n_32_585;
	 wire n_32_586;
	 wire n_32_587;
	 wire n_32_588;
	 wire n_32_589;
	 wire n_32_590;
	 wire n_32_591;
	 wire n_32_592;
	 wire n_32_593;
	 wire n_32_594;
	 wire n_32_595;
	 wire n_32_596;
	 wire n_32_597;
	 wire n_32_598;
	 wire n_32_599;
	 wire n_32_600;
	 wire n_32_601;
	 wire n_32_602;
	 wire n_32_603;
	 wire n_32_604;
	 wire n_32_605;
	 wire n_32_606;
	 wire n_32_607;
	 wire n_32_608;
	 wire n_32_609;
	 wire n_32_610;
	 wire n_32_611;
	 wire n_32_612;
	 wire n_32_613;
	 wire n_32_614;
	 wire n_32_615;
	 wire n_32_616;
	 wire n_32_617;
	 wire n_32_618;
	 wire n_32_619;
	 wire n_32_620;
	 wire n_32_621;
	 wire n_32_622;
	 wire n_32_623;
	 wire n_32_624;
	 wire n_32_625;
	 wire n_32_626;
	 wire n_32_627;
	 wire n_32_628;
	 wire n_32_629;
	 wire n_32_630;
	 wire n_32_631;
	 wire n_32_632;
	 wire n_32_633;
	 wire n_32_634;
	 wire n_32_635;
	 wire n_32_636;
	 wire n_32_637;
	 wire n_32_638;
	 wire n_32_639;
	 wire n_32_640;
	 wire n_32_641;
	 wire n_32_642;
	 wire n_32_643;
	 wire n_32_644;
	 wire n_32_645;
	 wire n_32_646;
	 wire n_32_647;
	 wire n_32_648;
	 wire n_32_649;
	 wire n_32_650;
	 wire n_32_651;
	 wire n_32_652;
	 wire n_32_653;
	 wire n_32_654;
	 wire n_32_655;
	 wire n_32_656;
	 wire n_32_657;
	 wire n_32_658;
	 wire n_32_659;
	 wire n_32_660;
	 wire n_32_661;
	 wire n_32_662;
	 wire n_32_663;
	 wire n_32_664;
	 wire n_32_665;
	 wire n_32_666;
	 wire n_32_667;
	 wire n_32_668;
	 wire n_32_669;
	 wire n_32_670;
	 wire n_32_671;
	 wire n_32_672;
	 wire n_32_673;
	 wire n_32_674;
	 wire n_34_0;
	 wire [31:0]product_xp;
	 wire n_34_1;
	 wire n_34_2;
	 wire n_34_3;
	 wire n_34_4;
	 wire n_34_5;
	 wire n_34_6;
	 wire n_34_7;
	 wire n_34_8;
	 wire n_34_9;
	 wire n_34_10;
	 wire n_34_11;
	 wire n_34_12;
	 wire n_34_13;
	 wire n_34_14;
	 wire n_34_15;
	 wire n_34_16;
	 wire n_34_17;
	 wire n_34_18;
	 wire n_34_19;
	 wire n_34_20;
	 wire n_34_21;
	 wire n_34_22;
	 wire n_34_23;
	 wire n_34_24;
	 wire n_34_25;
	 wire acc_sel;
	 wire n_38_0;
	 wire result_clr;
	 wire n_39_0;
	 wire n_39_1;
	 wire [15:0]reshi;
	 wire n_41_0;
	 wire n_41_1;
	 wire n_41_2;
	 wire n_41_3;
	 wire n_41_4;
	 wire n_41_5;
	 wire n_41_6;
	 wire n_41_7;
	 wire n_41_8;
	 wire n_41_9;
	 wire n_41_10;
	 wire n_41_11;
	 wire n_41_12;
	 wire n_41_13;
	 wire n_41_14;
	 wire n_41_15;
	 wire n_41_16;
	 wire n_42_0;
	 wire n_42_1;
	 wire n_45_0;
	 wire n_45_1;
	 wire n_45_2;
	 wire n_45_3;
	 wire n_45_4;
	 wire n_45_5;
	 wire n_45_6;
	 wire n_45_7;
	 wire n_45_8;
	 wire n_45_9;
	 wire n_45_10;
	 wire n_45_11;
	 wire n_45_12;
	 wire n_45_13;
	 wire n_45_14;
	 wire n_45_15;
	 wire n_45_16;
	 wire n_46_0;
	 wire n_46_1;
	 wire n_48_0;
	 wire n_48_1;
	 wire n_48_2;
	 wire n_48_3;
	 wire n_48_4;
	 wire n_48_5;
	 wire n_48_6;
	 wire n_48_7;
	 wire n_48_8;
	 wire n_48_9;
	 wire n_48_10;
	 wire n_48_11;
	 wire n_48_12;
	 wire n_48_13;
	 wire n_48_14;
	 wire n_48_15;
	 wire [15:0]reshi_nxt;
	 wire n_48_16;
	 wire n_48_17;
	 wire n_48_18;
	 wire n_48_19;
	 wire n_48_20;
	 wire n_48_21;
	 wire n_48_22;
	 wire n_48_23;
	 wire n_48_24;
	 wire n_48_25;
	 wire n_48_26;
	 wire n_48_27;
	 wire n_48_28;
	 wire n_48_29;
	 wire n_48_30;
	 wire n_50_0;
	 wire n_50_1;
	 wire [1:0]sumext_s_nxt;
	 wire [1:0]sumext_s;
	 wire n_52_0;
	 wire n_53_0;
	 wire n_53_1;
	 wire n_55_0;
	 wire n_55_1;
	 wire n_55_2;
	 wire n_57_0;
	 wire n_57_1;
	 wire n_60_0;
	 wire n_60_1;
	 wire n_60_2;
	 wire n_60_3;
	 wire n_60_4;
	 wire n_60_5;
	 wire n_60_6;
	 wire n_60_7;
	 wire n_60_8;
	 wire n_60_9;
	 wire n_60_10;
	 wire n_60_11;
	 wire n_60_12;
	 wire n_60_13;
	 wire n_60_14;
	 wire n_60_15;
	 wire n_60_16;
	 wire n_60_17;
	 wire n_60_18;
	 wire n_60_19;
	 wire n_60_20;
	 wire n_60_21;
	 wire n_60_22;
	 wire n_60_23;
	 wire n_60_24;
	 wire n_60_25;
	 wire n_60_26;
	 wire n_60_27;
	 wire n_60_28;
	 wire n_60_29;
	 wire n_60_30;
	 wire n_60_31;
	 wire n_60_32;
	 wire n_60_33;
	 wire n_60_34;
	 wire n_60_35;
	 wire n_60_36;
	 wire n_60_37;
	 wire n_60_38;
	 wire n_60_39;
	 wire n_60_40;
	 wire n_60_41;
	 wire n_60_42;
	 wire n_60_43;
	 wire n_60_44;
	 wire n_60_45;
	 wire n_60_46;
	 wire n_60_47;
	 wire n_60_48;
	 wire n_60_49;
	 wire n_60_50;
	 wire n_60_51;
	 wire n_60_52;
	 wire n_60_53;
	 wire n_60_54;
	 wire n_60_55;
	 wire n_60_56;
	 wire n_60_57;
	 wire n_60_58;
	 wire n_60_59;
	 wire n_60_60;
	 wire n_60_61;
	 wire n_60_62;
	 wire n_60_63;
	 wire n_60_64;
	 wire n_60_65;
	 wire n_60_66;
	 wire n_60_67;
	 wire n_60_68;
	 wire n_60_69;
	 wire n_60_70;
	 wire n_60_71;
	 wire n_60_72;
	 wire n_60_73;
	 wire n_60_74;
	 wire n_60_75;
	 wire n_60_76;
	 wire n_60_77;
	 wire n_60_78;
	 wire n_60_79;
	 wire n_60_80;
	 wire n_60_81;
	 wire n_60_82;
	 wire n_15;
	 wire n_5;
	 wire n_38;
	 wire n_3;
	 wire n_18;
	 wire n_4;
	 wire n_19;
	 wire n_68;
	 wire n_1;
	 wire n_16;
	 wire n_2;
	 wire n_17;
	 wire n_67;
	 wire n_6;
	 wire n_20;
	 wire n_21;
	 wire n_41;
	 wire n_45;
	 wire n_46;
	 wire n_47;
	 wire n_48;
	 wire n_49;
	 wire n_40;
	 wire n_39;
	 wire n_50;
	 wire n_51;
	 wire n_52;
	 wire n_53;
	 wire n_54;
	 wire n_55;
	 wire n_56;
	 wire n_57;
	 wire n_136;
	 wire n_119;
	 wire n_69;
	 wire n_121;
	 wire n_88;
	 wire n_90;
	 wire n_135;
	 wire n_118;
	 wire n_91;
	 wire n_134;
	 wire n_117;
	 wire n_92;
	 wire n_133;
	 wire n_116;
	 wire n_93;
	 wire n_44;
	 wire n_132;
	 wire n_115;
	 wire n_94;
	 wire n_43;
	 wire n_131;
	 wire n_114;
	 wire n_95;
	 wire n_42;
	 wire n_130;
	 wire n_113;
	 wire n_96;
	 wire n_129;
	 wire n_112;
	 wire n_97;
	 wire n_128;
	 wire n_111;
	 wire n_98;
	 wire n_127;
	 wire n_110;
	 wire n_99;
	 wire n_126;
	 wire n_109;
	 wire n_100;
	 wire n_125;
	 wire n_108;
	 wire n_101;
	 wire n_124;
	 wire n_107;
	 wire n_102;
	 wire n_123;
	 wire n_106;
	 wire n_103;
	 wire n_122;
	 wire n_105;
	 wire n_104;
	 wire n_89;
	 wire n_137;
	 wire n_120;
	 wire n_0;
	 wire n_13;
	 wire n_9;
	 wire n_11;
	 wire n_10;
	 wire n_150;
	 wire n_58;
	 wire n_59;
	 wire n_60;
	 wire n_61;
	 wire n_62;
	 wire n_63;
	 wire n_64;
	 wire n_65;
	 wire n_66;
	 wire n_7;
	 wire n_86;
	 wire n_87;
	 wire n_70;
	 wire n_85;
	 wire n_84;
	 wire n_83;
	 wire n_82;
	 wire n_81;
	 wire n_80;
	 wire n_79;
	 wire n_78;
	 wire n_77;
	 wire n_76;
	 wire n_75;
	 wire n_74;
	 wire n_73;
	 wire n_72;
	 wire n_71;
	 wire n_138;
	 wire n_142;
	 wire n_143;
	 wire n_140;
	 wire n_148;
	 wire n_8;
	 wire n_149;
	 wire n_12;
	 wire n_37;
	 wire n_14;
	 wire n_36;
	 wire n_35;
	 wire n_34;
	 wire n_33;
	 wire n_32;
	 wire n_31;
	 wire n_30;
	 wire n_29;
	 wire n_28;
	 wire n_27;
	 wire n_26;
	 wire n_25;
	 wire n_24;
	 wire n_145;
	 wire n_147;
	 wire n_23;
	 wire n_139;
	 wire n_141;
	 wire n_144;
	 wire n_146;
	 wire n_22;

endmodule

module omsp_and_gate__1_3(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_dbg_uart(dbg_addr,dbg_din,dbg_rd,dbg_uart_txd,dbg_wr,dbg_clk,dbg_dout,dbg_rd_rdy,dbg_rst,dbg_uart_rxd,mem_burst,mem_burst_end,mem_burst_rd,mem_burst_wr,mem_bw);
	 output [5:0]dbg_addr;
	 output [15:0]dbg_din;
	 output dbg_rd;
	 output dbg_uart_txd;
	 output dbg_wr;
	 input dbg_clk;
	 input [15:0]dbg_dout;
	 input dbg_rd_rdy;
	 input dbg_rst;
	 input dbg_uart_rxd;
	 input mem_burst;
	 input mem_burst_end;
	 input mem_burst_rd;
	 input mem_burst_wr;
	 input mem_bw;

	 wire uart_rxd_n;
	 wire uart_rxd;
	 wire [1:0]rxd_buf;
	 wire n_2_0;
	 wire n_2_1;
	 wire n_2_2;
	 wire rxd_maj_nxt;
	 wire [19:0]xfer_buf;
	 wire n_4_0;
	 wire n_4_1;
	 wire n_4_2;
	 wire n_4_3;
	 wire n_4_4;
	 wire n_4_5;
	 wire n_4_6;
	 wire n_4_7;
	 wire n_4_8;
	 wire n_4_9;
	 wire n_4_10;
	 wire n_4_11;
	 wire n_4_12;
	 wire n_4_13;
	 wire n_4_14;
	 wire n_4_15;
	 wire n_4_16;
	 wire n_4_17;
	 wire n_4_18;
	 wire n_5_0;
	 wire n_5_1;
	 wire rxd_maj;
	 wire n_7_0;
	 wire n_8_0;
	 wire n_8_1;
	 wire n_8_2;
	 wire n_8_3;
	 wire n_8_4;
	 wire n_8_5;
	 wire n_8_6;
	 wire n_8_7;
	 wire n_8_8;
	 wire n_8_9;
	 wire n_8_10;
	 wire n_8_11;
	 wire n_8_12;
	 wire n_8_13;
	 wire n_8_14;
	 wire n_8_15;
	 wire n_8_16;
	 wire n_8_17;
	 wire n_8_18;
	 wire n_8_19;
	 wire n_8_20;
	 wire n_8_21;
	 wire n_8_22;
	 wire n_8_23;
	 wire n_8_24;
	 wire [2:0]uart_state_nxt_reg;
	 wire n_8_25;
	 wire n_8_26;
	 wire n_8_27;
	 wire n_8_28;
	 wire n_8_29;
	 wire [2:0]uart_state;
	 wire n_11_0;
	 wire n_11_1;
	 wire n_13_0;
	 wire n_13_1;
	 wire n_13_2;
	 wire n_14_0;
	 wire n_15_0;
	 wire rxd_fe;
	 wire sync_busy;
	 wire [15:0]bit_cnt_max;
	 wire n_21_0;
	 wire n_21_1;
	 wire n_21_2;
	 wire n_21_3;
	 wire n_21_4;
	 wire n_21_5;
	 wire n_21_6;
	 wire n_21_7;
	 wire n_21_8;
	 wire n_21_9;
	 wire n_21_10;
	 wire n_21_11;
	 wire n_21_12;
	 wire n_21_13;
	 wire n_21_14;
	 wire n_21_15;
	 wire n_21_16;
	 wire n_21_17;
	 wire n_22_0;
	 wire n_22_1;
	 wire n_24_0;
	 wire txd_start;
	 wire rx_active;
	 wire [15:0]xfer_cnt;
	 wire n_27_0;
	 wire n_27_1;
	 wire n_27_2;
	 wire n_27_3;
	 wire n_27_4;
	 wire n_27_5;
	 wire n_27_6;
	 wire n_27_7;
	 wire n_27_8;
	 wire n_27_9;
	 wire n_27_10;
	 wire n_27_11;
	 wire n_27_12;
	 wire n_27_13;
	 wire n_29_0;
	 wire n_30_0;
	 wire n_31_0;
	 wire n_31_1;
	 wire n_31_2;
	 wire n_31_3;
	 wire n_31_4;
	 wire n_31_5;
	 wire n_31_6;
	 wire n_31_7;
	 wire n_31_8;
	 wire n_31_9;
	 wire n_31_10;
	 wire n_31_11;
	 wire n_31_12;
	 wire n_31_13;
	 wire n_31_14;
	 wire n_31_15;
	 wire n_31_16;
	 wire n_31_17;
	 wire n_31_18;
	 wire n_31_19;
	 wire n_31_20;
	 wire n_31_21;
	 wire n_31_22;
	 wire n_31_23;
	 wire n_31_24;
	 wire n_31_25;
	 wire n_31_26;
	 wire n_31_27;
	 wire n_31_28;
	 wire n_31_29;
	 wire n_31_30;
	 wire n_31_31;
	 wire n_31_32;
	 wire n_32_0;
	 wire n_32_1;
	 wire n_32_2;
	 wire n_32_3;
	 wire n_33_0;
	 wire n_33_1;
	 wire n_33_2;
	 wire n_35_0;
	 wire n_35_1;
	 wire n_35_2;
	 wire n_35_3;
	 wire n_35_4;
	 wire n_35_5;
	 wire xfer_bit_inc;
	 wire [3:0]xfer_bit;
	 wire n_39_0;
	 wire n_39_1;
	 wire n_39_2;
	 wire n_40_0;
	 wire n_41_0;
	 wire n_41_1;
	 wire n_42_0;
	 wire n_42_1;
	 wire n_42_2;
	 wire n_44_0;
	 wire n_44_1;
	 wire n_44_2;
	 wire n_44_3;
	 wire xfer_done;
	 wire cmd_valid;
	 wire dbg_bw;
	 wire n_49_0;
	 wire n_49_1;
	 wire n_49_2;
	 wire n_49_3;
	 wire n_49_4;
	 wire n_49_5;
	 wire n_49_6;
	 wire n_49_7;
	 wire n_49_8;
	 wire n_49_9;
	 wire n_49_10;
	 wire n_50_0;
	 wire n_50_1;
	 wire n_52_0;
	 wire n_52_1;
	 wire n_54_0;
	 wire n_136;
	 wire n_130;
	 wire n_19;
	 wire n_76;
	 wire n_53;
	 wire n_58;
	 wire n_54;
	 wire n_56;
	 wire n_57;
	 wire n_55;
	 wire n_52;
	 wire n_59;
	 wire n_51;
	 wire n_22;
	 wire n_119;
	 wire n_123;
	 wire n_124;
	 wire n_128;
	 wire n_118;
	 wire n_120;
	 wire n_125;
	 wire n_121;
	 wire n_122;
	 wire n_127;
	 wire n_116;
	 wire n_117;
	 wire n_28;
	 wire n_126;
	 wire n_25;
	 wire n_27;
	 wire n_26;
	 wire n_29;
	 wire n_31;
	 wire n_24;
	 wire n_23;
	 wire n_33;
	 wire n_34;
	 wire n_32;
	 wire n_50;
	 wire n_60;
	 wire n_61;
	 wire n_49;
	 wire n_95;
	 wire n_94;
	 wire n_97;
	 wire n_78;
	 wire n_96;
	 wire n_98;
	 wire n_79;
	 wire n_62;
	 wire n_48;
	 wire n_99;
	 wire n_77;
	 wire n_80;
	 wire n_63;
	 wire n_47;
	 wire n_100;
	 wire n_81;
	 wire n_64;
	 wire n_46;
	 wire n_101;
	 wire n_82;
	 wire n_65;
	 wire n_45;
	 wire n_102;
	 wire n_83;
	 wire n_66;
	 wire n_44;
	 wire n_103;
	 wire n_84;
	 wire n_67;
	 wire n_43;
	 wire n_104;
	 wire n_85;
	 wire n_68;
	 wire n_42;
	 wire n_105;
	 wire n_86;
	 wire n_69;
	 wire n_41;
	 wire n_106;
	 wire n_87;
	 wire n_70;
	 wire n_40;
	 wire n_107;
	 wire n_88;
	 wire n_71;
	 wire n_39;
	 wire n_108;
	 wire n_89;
	 wire n_72;
	 wire n_38;
	 wire n_109;
	 wire n_90;
	 wire n_73;
	 wire n_37;
	 wire n_110;
	 wire n_91;
	 wire n_74;
	 wire n_36;
	 wire n_111;
	 wire n_92;
	 wire n_75;
	 wire n_35;
	 wire n_112;
	 wire n_93;
	 wire n_113;
	 wire n_114;
	 wire n_115;
	 wire n_21;
	 wire n_0;
	 wire n_18;
	 wire n_17;
	 wire n_129;
	 wire n_16;
	 wire n_15;
	 wire n_14;
	 wire n_13;
	 wire n_12;
	 wire n_131;
	 wire n_11;
	 wire n_10;
	 wire n_20;
	 wire n_9;
	 wire n_8;
	 wire n_7;
	 wire n_6;
	 wire n_5;
	 wire n_4;
	 wire n_132;
	 wire n_30;
	 wire n_133;
	 wire n_3;
	 wire n_2;
	 wire n_1;
	 wire n_135;
	 wire n_134;

endmodule

module omsp_frontend(cpu_halt_st,decode_noirq,e_state,exec_done,inst_ad,inst_as,inst_alu,inst_bw,inst_dest,inst_dext,inst_irq_rst,inst_jmp,inst_mov,inst_sext,inst_so,inst_src,inst_type,irq_acc,mab,mb_en,mclk_dma_enable,mclk_dma_wkup,mclk_enable,mclk_wkup,nmi_acc,pc,pc_nxt,cpu_en_s,cpu_halt_cmd,cpuoff,dbg_reg_sel,dma_en,dma_wkup,fe_pmem_wait,gie,irq,mclk,mdb_in,nmi_pnd,nmi_wkup,pc_sw,pc_sw_wr,puc_rst,scan_enable,wdt_irq,wdt_wkup,wkup);
	 output cpu_halt_st;
	 output decode_noirq;
	 output [3:0]e_state;
	 output exec_done;
	 output [7:0]inst_ad;
	 output [7:0]inst_as;
	 output [11:0]inst_alu;
	 output inst_bw;
	 output [15:0]inst_dest;
	 output [15:0]inst_dext;
	 output inst_irq_rst;
	 output [7:0]inst_jmp;
	 output inst_mov;
	 output [15:0]inst_sext;
	 output [7:0]inst_so;
	 output [15:0]inst_src;
	 output [2:0]inst_type;
	 output [13:0]irq_acc;
	 output [15:0]mab;
	 output mb_en;
	 output mclk_dma_enable;
	 output mclk_dma_wkup;
	 output mclk_enable;
	 output mclk_wkup;
	 output nmi_acc;
	 output [15:0]pc;
	 output [15:0]pc_nxt;
	 input cpu_en_s;
	 input cpu_halt_cmd;
	 input cpuoff;
	 input [3:0]dbg_reg_sel;
	 input dma_en;
	 input dma_wkup;
	 input fe_pmem_wait;
	 input gie;
	 input [13:0]irq;
	 input mclk;
	 input [15:0]mdb_in;
	 input nmi_pnd;
	 input nmi_wkup;
	 input [15:0]pc_sw;
	 input pc_sw_wr;
	 input puc_rst;
	 input scan_enable;
	 input wdt_irq;
	 input wdt_wkup;
	 input wkup;

	 wire mirq_wkup;
	 wire n_0_0;
	 wire cpu_halt_req;
	 wire n_3_0;
	 wire n_3_1;
	 wire n_3_2;
	 wire n_3_3;
	 wire n_4_0;
	 wire n_4_1;
	 wire n_4_2;
	 wire [2:0]i_state;
	 wire n_6_0;
	 wire n_6_1;
	 wire n_6_2;
	 wire n_10_0;
	 wire n_10_1;
	 wire [3:0]src_reg;
	 wire n_10_2;
	 wire n_10_3;
	 wire n_10_4;
	 wire n_11_0;
	 wire inst_type_nxt;
	 wire n_12_0;
	 wire n_12_1;
	 wire n_12_2;
	 wire n_12_3;
	 wire n_12_4;
	 wire n_12_5;
	 wire n_12_6;
	 wire n_12_7;
	 wire n_12_8;
	 wire n_12_9;
	 wire [12:0]inst_as_nxt;
	 wire n_12_10;
	 wire n_12_11;
	 wire n_12_12;
	 wire n_12_13;
	 wire n_12_14;
	 wire n_13_0;
	 wire n_13_1;
	 wire is_const;
	 wire is_sext;
	 wire n_16_0;
	 wire inst_dext_rdy;
	 wire exec_dext_rdy;
	 wire n_19_0;
	 wire n_19_1;
	 wire n_20_0;
	 wire n_20_1;
	 wire n_20_2;
	 wire n_20_3;
	 wire n_22_0;
	 wire n_23_0;
	 wire n_23_1;
	 wire n_23_2;
	 wire n_23_3;
	 wire n_23_4;
	 wire n_23_5;
	 wire n_23_6;
	 wire n_23_7;
	 wire n_23_8;
	 wire n_23_9;
	 wire n_23_10;
	 wire n_23_11;
	 wire n_23_12;
	 wire n_23_13;
	 wire n_23_14;
	 wire n_23_15;
	 wire n_23_16;
	 wire n_23_17;
	 wire inst_ad_nxt;
	 wire n_25_0;
	 wire n_25_1;
	 wire n_25_2;
	 wire n_25_3;
	 wire n_25_4;
	 wire n_25_5;
	 wire n_25_6;
	 wire n_27_0;
	 wire [7:0]inst_so_nxt;
	 wire n_27_1;
	 wire inst_sext_rdy;
	 wire exec_dst_wr;
	 wire n_32_0;
	 wire n_33_0;
	 wire n_33_1;
	 wire n_33_2;
	 wire n_33_3;
	 wire n_33_4;
	 wire exec_src_wr;
	 wire n_39_0;
	 wire n_39_1;
	 wire exec_jmp;
	 wire n_44_0;
	 wire n_44_1;
	 wire n_45_0;
	 wire n_45_1;
	 wire n_45_2;
	 wire dst_acalc_pre;
	 wire src_acalc_pre;
	 wire n_50_0;
	 wire n_50_1;
	 wire n_50_2;
	 wire n_50_3;
	 wire n_50_4;
	 wire n_50_5;
	 wire n_50_6;
	 wire n_50_7;
	 wire n_50_8;
	 wire n_50_9;
	 wire n_50_10;
	 wire n_50_11;
	 wire n_50_12;
	 wire n_50_13;
	 wire n_50_14;
	 wire n_50_15;
	 wire n_50_16;
	 wire n_50_17;
	 wire n_50_18;
	 wire n_50_19;
	 wire n_53_0;
	 wire n_53_1;
	 wire n_55_0;
	 wire n_55_1;
	 wire n_55_2;
	 wire n_55_3;
	 wire n_55_4;
	 wire n_55_5;
	 wire n_55_6;
	 wire n_55_7;
	 wire n_55_8;
	 wire n_55_9;
	 wire n_55_10;
	 wire n_55_11;
	 wire n_55_12;
	 wire n_55_13;
	 wire n_55_14;
	 wire n_55_15;
	 wire n_55_16;
	 wire n_55_17;
	 wire n_55_18;
	 wire n_55_19;
	 wire n_55_20;
	 wire n_55_21;
	 wire n_55_22;
	 wire n_55_23;
	 wire n_55_24;
	 wire n_55_25;
	 wire n_55_26;
	 wire n_55_27;
	 wire n_55_28;
	 wire n_55_29;
	 wire n_55_30;
	 wire n_55_31;
	 wire n_55_32;
	 wire n_55_33;
	 wire n_55_34;
	 wire [3:0]e_state_nxt_reg;
	 wire n_55_35;
	 wire n_55_36;
	 wire n_55_37;
	 wire n_55_38;
	 wire n_55_39;
	 wire n_55_40;
	 wire n_55_41;
	 wire n_55_42;
	 wire n_55_43;
	 wire n_55_44;
	 wire n_55_45;
	 wire n_55_46;
	 wire n_55_47;
	 wire n_55_48;
	 wire n_55_49;
	 wire n_55_50;
	 wire n_55_51;
	 wire n_55_52;
	 wire n_55_53;
	 wire n_55_54;
	 wire n_55_55;
	 wire n_55_56;
	 wire n_55_57;
	 wire n_55_58;
	 wire n_55_59;
	 wire n_55_60;
	 wire n_55_61;
	 wire n_55_62;
	 wire n_55_63;
	 wire n_55_64;
	 wire n_55_65;
	 wire n_55_66;
	 wire n_55_67;
	 wire n_55_68;
	 wire n_58_0;
	 wire n_58_1;
	 wire n_58_2;
	 wire n_58_3;
	 wire n_59_0;
	 wire n_59_1;
	 wire n_59_2;
	 wire n_59_3;
	 wire n_59_4;
	 wire n_59_5;
	 wire n_59_6;
	 wire n_60_0;
	 wire irq_detect;
	 wire decode;
	 wire n_64_0;
	 wire [1:0]inst_sz_nxt;
	 wire [1:0]inst_sz;
	 wire n_70_0;
	 wire n_71_0;
	 wire n_72_0;
	 wire n_73_0;
	 wire n_73_1;
	 wire n_73_2;
	 wire n_73_3;
	 wire n_74_0;
	 wire n_75_0;
	 wire n_76_0;
	 wire n_76_1;
	 wire n_76_2;
	 wire n_76_3;
	 wire n_76_4;
	 wire n_76_5;
	 wire n_76_6;
	 wire n_76_7;
	 wire [2:0]i_state_nxt_reg;
	 wire n_76_8;
	 wire n_76_9;
	 wire n_76_10;
	 wire n_76_11;
	 wire n_76_12;
	 wire n_76_13;
	 wire n_76_14;
	 wire n_80_0;
	 wire n_82_0;
	 wire n_82_1;
	 wire n_82_2;
	 wire n_82_3;
	 wire n_82_4;
	 wire n_82_5;
	 wire n_82_6;
	 wire n_82_7;
	 wire n_82_8;
	 wire n_82_9;
	 wire n_82_10;
	 wire [11:0]inst_to_nxt;
	 wire alu_inc;
	 wire [11:0]inst_alu_nxt;
	 wire n_88_0;
	 wire n_88_1;
	 wire n_91_0;
	 wire [3:0]inst_dest_bin;
	 wire n_94_0;
	 wire n_94_1;
	 wire n_94_2;
	 wire n_94_3;
	 wire n_94_4;
	 wire n_94_5;
	 wire n_94_6;
	 wire n_94_7;
	 wire n_94_8;
	 wire n_94_9;
	 wire n_94_10;
	 wire n_94_11;
	 wire n_95_0;
	 wire n_95_1;
	 wire n_95_2;
	 wire n_95_3;
	 wire n_95_4;
	 wire n_95_5;
	 wire n_95_6;
	 wire n_95_7;
	 wire n_95_8;
	 wire n_95_9;
	 wire n_95_10;
	 wire n_95_11;
	 wire n_97_0;
	 wire n_97_1;
	 wire n_97_2;
	 wire n_97_3;
	 wire n_97_4;
	 wire n_97_5;
	 wire n_97_6;
	 wire n_97_7;
	 wire n_97_8;
	 wire n_97_9;
	 wire n_97_10;
	 wire n_97_11;
	 wire n_97_12;
	 wire n_97_13;
	 wire n_97_14;
	 wire n_97_15;
	 wire n_97_16;
	 wire n_97_17;
	 wire n_97_18;
	 wire n_97_19;
	 wire n_98_0;
	 wire n_98_1;
	 wire n_98_2;
	 wire n_98_3;
	 wire n_98_4;
	 wire n_99_0;
	 wire [15:0]ext_nxt;
	 wire n_99_1;
	 wire n_99_2;
	 wire n_99_3;
	 wire n_99_4;
	 wire n_99_5;
	 wire n_99_6;
	 wire n_99_7;
	 wire n_99_8;
	 wire n_99_9;
	 wire n_99_10;
	 wire n_99_11;
	 wire n_99_12;
	 wire n_99_13;
	 wire n_99_14;
	 wire n_99_15;
	 wire n_99_16;
	 wire n_99_17;
	 wire n_101_0;
	 wire n_101_1;
	 wire [2:0]inst_jmp_bin;
	 wire n_105_0;
	 wire n_105_1;
	 wire n_105_2;
	 wire n_105_3;
	 wire n_105_4;
	 wire n_105_5;
	 wire n_105_6;
	 wire n_110_0;
	 wire n_110_1;
	 wire n_110_2;
	 wire n_110_3;
	 wire n_110_4;
	 wire n_110_5;
	 wire n_110_6;
	 wire n_110_7;
	 wire n_110_8;
	 wire n_110_9;
	 wire n_110_10;
	 wire n_110_11;
	 wire n_110_12;
	 wire n_110_13;
	 wire n_110_14;
	 wire n_110_15;
	 wire n_110_16;
	 wire n_110_17;
	 wire n_110_18;
	 wire n_110_19;
	 wire n_110_20;
	 wire n_110_21;
	 wire n_110_22;
	 wire n_110_23;
	 wire n_110_24;
	 wire n_110_25;
	 wire n_110_26;
	 wire n_110_27;
	 wire n_110_28;
	 wire n_110_29;
	 wire n_110_30;
	 wire n_110_31;
	 wire n_110_32;
	 wire n_110_33;
	 wire n_110_34;
	 wire n_110_35;
	 wire n_111_0;
	 wire n_111_1;
	 wire n_111_2;
	 wire n_111_3;
	 wire n_111_4;
	 wire [3:0]inst_src_bin;
	 wire n_114_0;
	 wire n_114_1;
	 wire n_114_2;
	 wire n_114_3;
	 wire n_114_4;
	 wire n_114_5;
	 wire n_114_6;
	 wire n_114_7;
	 wire n_114_8;
	 wire n_114_9;
	 wire n_114_10;
	 wire n_114_11;
	 wire n_115_0;
	 wire n_115_1;
	 wire n_115_2;
	 wire n_115_3;
	 wire n_115_4;
	 wire n_115_5;
	 wire n_115_6;
	 wire n_115_7;
	 wire n_115_8;
	 wire n_115_9;
	 wire n_115_10;
	 wire n_115_11;
	 wire n_115_12;
	 wire n_115_13;
	 wire n_115_14;
	 wire n_115_15;
	 wire n_115_16;
	 wire n_115_17;
	 wire n_115_18;
	 wire n_115_19;
	 wire [5:0]irq_num;
	 wire n_118_0;
	 wire n_118_1;
	 wire n_118_2;
	 wire n_118_3;
	 wire n_118_4;
	 wire n_118_5;
	 wire n_118_6;
	 wire n_118_7;
	 wire n_118_8;
	 wire n_118_9;
	 wire n_118_10;
	 wire n_118_11;
	 wire n_118_12;
	 wire n_118_13;
	 wire n_118_14;
	 wire n_118_15;
	 wire n_118_16;
	 wire n_118_17;
	 wire n_118_18;
	 wire n_118_19;
	 wire n_118_20;
	 wire n_118_21;
	 wire n_118_22;
	 wire n_118_23;
	 wire n_118_24;
	 wire n_118_25;
	 wire n_118_26;
	 wire n_118_27;
	 wire n_118_28;
	 wire n_118_29;
	 wire n_118_30;
	 wire n_118_31;
	 wire n_118_32;
	 wire n_118_33;
	 wire n_118_34;
	 wire n_118_35;
	 wire n_118_36;
	 wire n_118_37;
	 wire n_118_38;
	 wire n_118_39;
	 wire n_118_40;
	 wire n_118_41;
	 wire n_118_42;
	 wire n_118_43;
	 wire n_118_44;
	 wire n_118_45;
	 wire n_118_46;
	 wire n_118_47;
	 wire n_118_48;
	 wire n_118_49;
	 wire n_118_50;
	 wire n_118_51;
	 wire n_118_52;
	 wire n_118_53;
	 wire n_118_54;
	 wire n_118_55;
	 wire n_118_56;
	 wire n_120_0;
	 wire n_120_1;
	 wire n_120_2;
	 wire n_120_3;
	 wire n_120_4;
	 wire n_120_5;
	 wire n_120_6;
	 wire n_120_7;
	 wire n_120_8;
	 wire n_120_9;
	 wire n_120_10;
	 wire n_120_11;
	 wire n_120_12;
	 wire n_120_13;
	 wire n_120_14;
	 wire n_120_15;
	 wire n_120_16;
	 wire n_120_17;
	 wire n_120_18;
	 wire n_120_19;
	 wire n_120_20;
	 wire n_122_0;
	 wire n_122_1;
	 wire n_122_2;
	 wire fetch;
	 wire [15:0]pc_incr;
	 wire n_124_0;
	 wire n_124_1;
	 wire n_124_2;
	 wire n_124_3;
	 wire n_124_4;
	 wire n_124_5;
	 wire n_124_6;
	 wire n_124_7;
	 wire n_124_8;
	 wire n_124_9;
	 wire n_124_10;
	 wire n_124_11;
	 wire n_124_12;
	 wire n_124_13;
	 wire n_124_14;
	 wire n_125_0;
	 wire n_126_0;
	 wire n_126_1;
	 wire n_126_2;
	 wire n_126_3;
	 wire n_126_4;
	 wire n_126_5;
	 wire n_126_6;
	 wire n_126_7;
	 wire n_126_8;
	 wire n_126_9;
	 wire n_126_10;
	 wire n_126_11;
	 wire n_126_12;
	 wire n_126_13;
	 wire n_126_14;
	 wire n_126_15;
	 wire n_127_0;
	 wire n_127_1;
	 wire n_127_2;
	 wire n_127_3;
	 wire n_127_4;
	 wire n_127_5;
	 wire n_127_6;
	 wire n_127_7;
	 wire n_127_8;
	 wire n_127_9;
	 wire n_127_10;
	 wire n_127_11;
	 wire n_127_12;
	 wire n_127_13;
	 wire n_127_14;
	 wire n_127_15;
	 wire n_127_16;
	 wire pmem_busy;
	 wire n_128_0;
	 wire n_128_1;
	 wire n_130_0;
	 wire n_130_1;
	 wire n_130_2;
	 wire n_130_3;
	 wire n_91;
	 wire n_0;
	 wire n_87;
	 wire n_1;
	 wire n_2;
	 wire n_3;
	 wire n_88;
	 wire n_89;
	 wire n_5;
	 wire n_55;
	 wire n_10;
	 wire n_29;
	 wire n_37;
	 wire n_28;
	 wire n_36;
	 wire n_9;
	 wire n_49;
	 wire n_17;
	 wire n_18;
	 wire n_48;
	 wire n_4;
	 wire n_67;
	 wire n_73;
	 wire n_51;
	 wire n_52;
	 wire n_50;
	 wire n_11;
	 wire n_43;
	 wire n_68;
	 wire n_45;
	 wire n_69;
	 wire n_70;
	 wire n_46;
	 wire n_47;
	 wire n_44;
	 wire n_72;
	 wire n_71;
	 wire n_56;
	 wire n_54;
	 wire n_20;
	 wire n_19;
	 wire n_26;
	 wire n_34;
	 wire n_27;
	 wire n_35;
	 wire n_53;
	 wire n_58;
	 wire n_6;
	 wire n_12;
	 wire n_38;
	 wire n_39;
	 wire n_62;
	 wire n_21;
	 wire n_63;
	 wire n_64;
	 wire n_57;
	 wire n_13;
	 wire n_7;
	 wire n_15;
	 wire n_16;
	 wire n_14;
	 wire n_61;
	 wire n_66;
	 wire n_65;
	 wire n_41;
	 wire n_42;
	 wire n_40;
	 wire n_59;
	 wire n_60;
	 wire n_82;
	 wire n_83;
	 wire n_86;
	 wire n_74;
	 wire n_75;
	 wire n_76;
	 wire n_79;
	 wire n_80;
	 wire n_90;
	 wire n_85;
	 wire n_81;
	 wire n_77;
	 wire n_78;
	 wire n_84;
	 wire n_92;
	 wire n_98;
	 wire n_100;
	 wire n_108;
	 wire n_24;
	 wire n_32;
	 wire n_22;
	 wire n_30;
	 wire n_104;
	 wire n_107;
	 wire n_25;
	 wire n_33;
	 wire n_94;
	 wire n_97;
	 wire n_96;
	 wire n_95;
	 wire n_105;
	 wire n_106;
	 wire n_103;
	 wire n_99;
	 wire n_102;
	 wire n_101;
	 wire n_110;
	 wire n_109;
	 wire n_144;
	 wire n_111;
	 wire n_127;
	 wire n_143;
	 wire n_126;
	 wire n_142;
	 wire n_125;
	 wire n_141;
	 wire n_124;
	 wire n_140;
	 wire n_123;
	 wire n_139;
	 wire n_122;
	 wire n_138;
	 wire n_121;
	 wire n_137;
	 wire n_120;
	 wire n_136;
	 wire n_119;
	 wire n_135;
	 wire n_118;
	 wire n_134;
	 wire n_117;
	 wire n_133;
	 wire n_116;
	 wire n_132;
	 wire n_115;
	 wire n_131;
	 wire n_114;
	 wire n_130;
	 wire n_113;
	 wire n_129;
	 wire n_112;
	 wire n_128;
	 wire n_145;
	 wire n_147;
	 wire n_146;
	 wire n_148;
	 wire n_149;
	 wire n_157;
	 wire n_156;
	 wire n_155;
	 wire n_154;
	 wire n_153;
	 wire n_152;
	 wire n_151;
	 wire n_150;
	 wire n_93;
	 wire n_158;
	 wire n_179;
	 wire n_180;
	 wire n_163;
	 wire n_178;
	 wire n_177;
	 wire n_176;
	 wire n_175;
	 wire n_174;
	 wire n_173;
	 wire n_172;
	 wire n_171;
	 wire n_170;
	 wire n_169;
	 wire n_168;
	 wire n_162;
	 wire n_167;
	 wire n_161;
	 wire n_166;
	 wire n_160;
	 wire n_165;
	 wire n_159;
	 wire n_164;
	 wire n_23;
	 wire n_31;
	 wire n_181;
	 wire n_197;
	 wire n_196;
	 wire n_195;
	 wire n_194;
	 wire n_193;
	 wire n_192;
	 wire n_191;
	 wire n_190;
	 wire n_189;
	 wire n_188;
	 wire n_187;
	 wire n_186;
	 wire n_185;
	 wire n_184;
	 wire n_183;
	 wire n_182;
	 wire n_8;
	 wire n_198;
	 wire n_200;
	 wire n_199;
	 wire n_201;
	 wire n_202;
	 wire n_203;
	 wire n_204;
	 wire n_218;
	 wire n_217;
	 wire n_216;
	 wire n_215;
	 wire n_214;
	 wire n_213;
	 wire n_212;
	 wire n_211;
	 wire n_210;
	 wire n_209;
	 wire n_208;
	 wire n_207;
	 wire n_206;
	 wire n_205;
	 wire n_221;
	 wire n_220;
	 wire n_222;
	 wire n_237;
	 wire n_236;
	 wire n_235;
	 wire n_234;
	 wire n_233;
	 wire n_232;
	 wire n_231;
	 wire n_230;
	 wire n_229;
	 wire n_228;
	 wire n_227;
	 wire n_226;
	 wire n_225;
	 wire n_224;
	 wire n_238;
	 wire n_223;
	 wire n_240;
	 wire n_239;
	 wire n_219;

endmodule

module OR4_X1_LVT(ZN,A1,A2,A3,A4);
	 output ZN;
	 input A1;
	 input A2;
	 input A3;
	 input A4;


endmodule

module omsp_sync_cell__2_21(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_and_gate__2_55(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_sfr(cpu_id,nmi_pnd,nmi_wkup,per_dout,wdtie,wdtifg_sw_clr,wdtifg_sw_set,cpu_nr_inst,cpu_nr_total,mclk,nmi,nmi_acc,per_addr,per_din,per_en,per_we,puc_rst,scan_mode,wdtifg,wdtnmies);
	 output [31:0]cpu_id;
	 output nmi_pnd;
	 output nmi_wkup;
	 output [15:0]per_dout;
	 output wdtie;
	 output wdtifg_sw_clr;
	 output wdtifg_sw_set;
	 input [7:0]cpu_nr_inst;
	 input [7:0]cpu_nr_total;
	 input mclk;
	 input nmi;
	 input nmi_acc;
	 input [13:0]per_addr;
	 input [15:0]per_din;
	 input per_en;
	 input [1:0]per_we;
	 input puc_rst;
	 input scan_mode;
	 input wdtifg;
	 input wdtnmies;

	 wire nmi_capture;
	 wire nmi_s;
	 wire n_0_0;
	 wire n_0_1;
	 wire n_0_2;
	 wire n_0_3;
	 wire reg_sel;
	 wire reg_lo_write;
	 wire n_2_0;
	 wire n_2_1;
	 wire n_2_2;
	 wire n_2_3;
	 wire n_2_4;
	 wire n_2_5;
	 wire n_2_6;
	 wire ifg1_wr;
	 wire nmi_capture_rst;
	 wire n_4_0;
	 wire nmie;
	 wire n_7_0;
	 wire n_8_0;
	 wire n_8_1;
	 wire nmi_dly;
	 wire n_10_0;
	 wire nmi_edge;
	 wire nmiifg;
	 wire n_13_0;
	 wire n_13_1;
	 wire n_14_0;
	 wire n_14_1;
	 wire reg_read;
	 wire n_27_0;
	 wire n_28_0;
	 wire nmi_pol;
	 wire n_1;
	 wire n_6;
	 wire n_11;
	 wire n_12;
	 wire n_13;
	 wire n_10;
	 wire n_8;
	 wire n_0;
	 wire n_5;
	 wire n_9;
	 wire n_7;
	 wire n_31;
	 wire n_14;
	 wire n_4;
	 wire n_19;
	 wire n_3;
	 wire n_18;
	 wire n_25;
	 wire n_2;
	 wire n_17;
	 wire n_24;
	 wire n_15;
	 wire n_30;
	 wire n_16;
	 wire n_27;
	 wire n_23;
	 wire n_22;
	 wire n_21;
	 wire n_26;
	 wire n_20;
	 wire n_28;
	 wire n_29;

endmodule

module omsp_and_gate__2_43(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_dbg(dbg_cpu_reset,dbg_freeze,dbg_halt_cmd,dbg_i2c_sda_out,dbg_mem_addr,dbg_mem_dout,dbg_mem_en,dbg_mem_wr,dbg_reg_wr,dbg_uart_txd,cpu_en_s,cpu_id,cpu_nr_inst,cpu_nr_total,dbg_clk,dbg_en_s,dbg_halt_st,dbg_i2c_addr,dbg_i2c_broadcast,dbg_i2c_scl,dbg_i2c_sda_in,dbg_mem_din,dbg_reg_din,dbg_rst,dbg_uart_rxd,decode_noirq,eu_mab,eu_mb_en,eu_mb_wr,fe_mdb_in,pc,puc_pnd_set);
	 output dbg_cpu_reset;
	 output dbg_freeze;
	 output dbg_halt_cmd;
	 output dbg_i2c_sda_out;
	 output [15:0]dbg_mem_addr;
	 output [15:0]dbg_mem_dout;
	 output dbg_mem_en;
	 output [1:0]dbg_mem_wr;
	 output dbg_reg_wr;
	 output dbg_uart_txd;
	 input cpu_en_s;
	 input [31:0]cpu_id;
	 input [7:0]cpu_nr_inst;
	 input [7:0]cpu_nr_total;
	 input dbg_clk;
	 input dbg_en_s;
	 input dbg_halt_st;
	 input [6:0]dbg_i2c_addr;
	 input [6:0]dbg_i2c_broadcast;
	 input dbg_i2c_scl;
	 input dbg_i2c_sda_in;
	 input [15:0]dbg_mem_din;
	 input [15:0]dbg_reg_din;
	 input dbg_rst;
	 input dbg_uart_rxd;
	 input decode_noirq;
	 input [15:0]eu_mab;
	 input eu_mb_en;
	 input [1:0]eu_mb_wr;
	 input [15:0]fe_mdb_in;
	 input [15:0]pc;
	 input puc_pnd_set;

	 wire dbg_wr;
	 wire dbg_rd;
	 wire [15:0]dbg_din;
	 wire [5:0]dbg_addr;
	 wire n_0_0;
	 wire n_0_1;
	 wire n_0_2;
	 wire n_0_3;
	 wire mem_start;
	 wire [2:0]mem_ctl;
	 wire mem_burst_rd;
	 wire mem_startb;
	 wire n_6_0;
	 wire n_6_1;
	 wire n_8_0;
	 wire n_9_0;
	 wire n_9_1;
	 wire n_9_2;
	 wire n_9_3;
	 wire n_9_4;
	 wire n_9_5;
	 wire [1:0]mem_state_nxt_reg;
	 wire n_9_6;
	 wire [1:0]mem_state;
	 wire n_12_0;
	 wire mem_access;
	 wire n_16_0;
	 wire n_17_0;
	 wire n_17_1;
	 wire n_17_2;
	 wire n_17_3;
	 wire n_17_4;
	 wire n_17_5;
	 wire n_17_6;
	 wire n_19_0;
	 wire n_19_1;
	 wire n_19_2;
	 wire n_19_3;
	 wire n_19_4;
	 wire n_19_5;
	 wire n_19_6;
	 wire n_19_7;
	 wire n_19_8;
	 wire n_19_9;
	 wire n_19_10;
	 wire n_19_11;
	 wire n_19_12;
	 wire n_19_13;
	 wire n_19_14;
	 wire n_19_15;
	 wire n_20_0;
	 wire n_20_1;
	 wire n_20_2;
	 wire n_20_3;
	 wire n_20_4;
	 wire n_20_5;
	 wire n_20_6;
	 wire n_20_7;
	 wire n_20_8;
	 wire n_20_9;
	 wire n_20_10;
	 wire n_20_11;
	 wire n_20_12;
	 wire n_20_13;
	 wire n_20_14;
	 wire n_20_15;
	 wire n_20_16;
	 wire n_22_0;
	 wire dbg_reg_rd;
	 wire dbg_mem_rd;
	 wire dbg_mem_rd_dly;
	 wire dbg_rd_rdy;
	 wire n_32_0;
	 wire n_32_1;
	 wire n_34_0;
	 wire dbg_mem_acc;
	 wire n_35_0;
	 wire n_35_1;
	 wire n_37_0;
	 wire n_37_1;
	 wire n_37_2;
	 wire n_37_3;
	 wire n_37_4;
	 wire [15:0]mem_cnt;
	 wire n_39_0;
	 wire n_39_1;
	 wire n_39_2;
	 wire n_39_3;
	 wire n_39_4;
	 wire n_39_5;
	 wire n_39_6;
	 wire n_39_7;
	 wire n_39_8;
	 wire n_39_9;
	 wire n_39_10;
	 wire n_39_11;
	 wire n_39_12;
	 wire n_39_13;
	 wire n_39_14;
	 wire n_39_15;
	 wire n_39_16;
	 wire n_40_0;
	 wire n_40_1;
	 wire n_40_2;
	 wire n_40_3;
	 wire n_40_4;
	 wire n_40_5;
	 wire n_40_6;
	 wire n_40_7;
	 wire n_40_8;
	 wire n_40_9;
	 wire n_40_10;
	 wire n_40_11;
	 wire n_40_12;
	 wire n_40_13;
	 wire n_40_14;
	 wire n_40_15;
	 wire n_40_16;
	 wire n_42_0;
	 wire n_42_1;
	 wire n_42_2;
	 wire n_42_3;
	 wire mem_burst_start;
	 wire n_44_0;
	 wire mem_burst_end;
	 wire mem_burst;
	 wire n_46_0;
	 wire n_46_1;
	 wire n_48_0;
	 wire [5:0]dbg_addr_in;
	 wire n_48_1;
	 wire n_48_2;
	 wire n_49_0;
	 wire n_49_1;
	 wire n_49_2;
	 wire n_49_3;
	 wire n_49_4;
	 wire n_49_5;
	 wire n_49_6;
	 wire n_49_7;
	 wire n_49_8;
	 wire n_49_9;
	 wire n_49_10;
	 wire n_49_11;
	 wire n_49_12;
	 wire n_49_13;
	 wire n_49_14;
	 wire n_49_15;
	 wire n_49_16;
	 wire n_49_17;
	 wire n_49_18;
	 wire n_49_19;
	 wire n_49_20;
	 wire n_49_21;
	 wire cpu_ctl_wr;
	 wire mem_ctl_wr;
	 wire mem_data_wr;
	 wire [3:0]cpu_ctl;
	 wire n_53_0;
	 wire n_53_1;
	 wire n_54_0;
	 wire n_54_1;
	 wire n_54_2;
	 wire n_54_3;
	 wire n_54_4;
	 wire dbg_swbrk;
	 wire n_55_0;
	 wire n_55_1;
	 wire n_55_2;
	 wire n_55_3;
	 wire n_55_4;
	 wire n_55_5;
	 wire halt_flag_set;
	 wire n_57_0;
	 wire n_57_1;
	 wire n_57_2;
	 wire halt_flag_clr;
	 wire halt_flag;
	 wire n_59_0;
	 wire n_60_0;
	 wire n_60_1;
	 wire istep;
	 wire n_64_0;
	 wire n_64_1;
	 wire n_66_0;
	 wire n_68_0;
	 wire n_68_1;
	 wire n_68_2;
	 wire n_68_3;
	 wire n_68_4;
	 wire n_68_5;
	 wire n_68_6;
	 wire n_68_7;
	 wire n_68_8;
	 wire [15:0]mem_data;
	 wire n_70_0;
	 wire n_71_0;
	 wire n_71_1;
	 wire n_71_2;
	 wire n_71_3;
	 wire n_71_4;
	 wire n_71_5;
	 wire n_71_6;
	 wire n_71_7;
	 wire n_71_8;
	 wire n_71_9;
	 wire n_71_10;
	 wire n_71_11;
	 wire n_71_12;
	 wire n_71_13;
	 wire n_71_14;
	 wire n_71_15;
	 wire n_72_0;
	 wire n_72_1;
	 wire n_72_2;
	 wire n_74_0;
	 wire n_74_1;
	 wire n_74_2;
	 wire n_74_3;
	 wire n_74_4;
	 wire n_74_5;
	 wire n_74_6;
	 wire n_74_7;
	 wire n_74_8;
	 wire n_74_9;
	 wire n_74_10;
	 wire n_74_11;
	 wire n_74_12;
	 wire n_74_13;
	 wire n_74_14;
	 wire n_74_15;
	 wire n_74_16;
	 wire n_74_17;
	 wire n_74_18;
	 wire n_74_19;
	 wire [1:0]cpu_stat;
	 wire n_76_0;
	 wire n_76_1;
	 wire n_76_2;
	 wire n_76_3;
	 wire n_76_4;
	 wire n_76_5;
	 wire n_76_6;
	 wire n_78_0;
	 wire n_78_1;
	 wire n_78_2;
	 wire n_78_3;
	 wire n_78_4;
	 wire n_78_5;
	 wire n_78_6;
	 wire n_78_7;
	 wire [15:0]dbg_dout;
	 wire n_78_8;
	 wire n_78_9;
	 wire n_78_10;
	 wire n_78_11;
	 wire n_78_12;
	 wire n_78_13;
	 wire n_78_14;
	 wire n_78_15;
	 wire n_78_16;
	 wire n_78_17;
	 wire n_78_18;
	 wire n_78_19;
	 wire n_78_20;
	 wire n_78_21;
	 wire n_78_22;
	 wire n_78_23;
	 wire n_78_24;
	 wire n_78_25;
	 wire n_78_26;
	 wire n_78_27;
	 wire n_78_28;
	 wire n_78_29;
	 wire n_78_30;
	 wire n_78_31;
	 wire n_78_32;
	 wire n_78_33;
	 wire n_78_34;
	 wire n_78_35;
	 wire n_78_36;
	 wire n_78_37;
	 wire n_78_38;
	 wire n_78_39;
	 wire n_78_40;
	 wire n_78_41;
	 wire n_78_42;
	 wire n_78_43;
	 wire n_78_44;
	 wire n_78_45;
	 wire n_78_46;
	 wire n_78_47;
	 wire n_78_48;
	 wire n_78_49;
	 wire n_78_50;
	 wire n_78_51;
	 wire n_78_52;
	 wire n_78_53;
	 wire n_78_54;
	 wire n_78_55;
	 wire n_78_56;
	 wire n_78_57;
	 wire n_78_58;
	 wire n_78_59;
	 wire n_78_60;
	 wire n_78_61;
	 wire n_78_62;
	 wire n_78_63;
	 wire n_78_64;
	 wire n_78_65;
	 wire n_78_66;
	 wire n_78_67;
	 wire n_78_68;
	 wire n_78_69;
	 wire n_78_70;
	 wire n_78_71;
	 wire n_78_72;
	 wire n_78_73;
	 wire n_78_74;
	 wire n_78_75;
	 wire n_78_76;
	 wire n_78_77;
	 wire n_78_78;
	 wire n_78_79;
	 wire n_78_80;
	 wire n_78_81;
	 wire n_78_82;
	 wire n_78_83;
	 wire n_78_84;
	 wire n_78_85;
	 wire n_78_86;
	 wire n_78_87;
	 wire n_78_88;
	 wire n_78_89;
	 wire n_78_90;
	 wire n_78_91;
	 wire n_78_92;
	 wire n_78_93;
	 wire n_78_94;
	 wire n_78_95;
	 wire n_78_96;
	 wire n_78_97;
	 wire n_78_98;
	 wire n_78_99;
	 wire n_78_100;
	 wire n_78_101;
	 wire n_78_102;
	 wire n_78_103;
	 wire n_78_104;
	 wire n_78_105;
	 wire n_78_106;
	 wire n_78_107;
	 wire n_78_108;
	 wire n_78_109;
	 wire n_78_110;
	 wire n_78_111;
	 wire n_78_112;
	 wire n_78_113;
	 wire n_78_114;
	 wire n_78_115;
	 wire mem_burst_wr;
	 wire n_95;
	 wire n_1;
	 wire n_104;
	 wire n_98;
	 wire n_102;
	 wire n_55;
	 wire n_57;
	 wire n_73;
	 wire n_58;
	 wire n_74;
	 wire n_59;
	 wire n_75;
	 wire n_60;
	 wire n_76;
	 wire n_61;
	 wire n_77;
	 wire n_62;
	 wire n_78;
	 wire n_63;
	 wire n_79;
	 wire n_64;
	 wire n_80;
	 wire n_65;
	 wire n_81;
	 wire n_66;
	 wire n_82;
	 wire n_67;
	 wire n_83;
	 wire n_68;
	 wire n_84;
	 wire n_69;
	 wire n_85;
	 wire n_70;
	 wire n_86;
	 wire n_71;
	 wire n_87;
	 wire n_2;
	 wire n_3;
	 wire n_4;
	 wire n_0;
	 wire n_5;
	 wire n_6;
	 wire n_7;
	 wire n_47;
	 wire n_48;
	 wire n_96;
	 wire n_101;
	 wire n_10;
	 wire n_53;
	 wire n_11;
	 wire n_13;
	 wire n_29;
	 wire n_46;
	 wire n_45;
	 wire n_49;
	 wire n_51;
	 wire n_9;
	 wire n_50;
	 wire n_52;
	 wire n_54;
	 wire n_56;
	 wire n_72;
	 wire n_88;
	 wire n_90;
	 wire n_89;
	 wire n_27;
	 wire n_43;
	 wire n_26;
	 wire n_42;
	 wire n_25;
	 wire n_41;
	 wire n_24;
	 wire n_40;
	 wire n_23;
	 wire n_39;
	 wire n_22;
	 wire n_38;
	 wire n_21;
	 wire n_37;
	 wire n_20;
	 wire n_36;
	 wire n_19;
	 wire n_35;
	 wire n_18;
	 wire n_34;
	 wire n_17;
	 wire n_33;
	 wire n_16;
	 wire n_32;
	 wire n_15;
	 wire n_31;
	 wire n_12;
	 wire n_14;
	 wire n_30;
	 wire n_28;
	 wire n_44;
	 wire n_97;
	 wire n_136;
	 wire n_135;
	 wire n_115;
	 wire n_133;
	 wire n_152;
	 wire n_153;
	 wire n_134;
	 wire n_92;
	 wire n_91;
	 wire n_99;
	 wire n_132;
	 wire n_151;
	 wire n_131;
	 wire n_150;
	 wire n_130;
	 wire n_149;
	 wire n_129;
	 wire n_148;
	 wire n_128;
	 wire n_147;
	 wire n_127;
	 wire n_146;
	 wire n_126;
	 wire n_145;
	 wire n_116;
	 wire n_117;
	 wire n_125;
	 wire n_144;
	 wire n_124;
	 wire n_143;
	 wire n_93;
	 wire n_123;
	 wire n_142;
	 wire n_105;
	 wire n_122;
	 wire n_141;
	 wire n_106;
	 wire n_121;
	 wire n_140;
	 wire n_94;
	 wire n_107;
	 wire n_100;
	 wire n_155;
	 wire n_120;
	 wire n_139;
	 wire n_154;
	 wire n_119;
	 wire n_138;
	 wire n_118;
	 wire n_137;
	 wire n_103;
	 wire n_8;
	 wire n_108;
	 wire n_110;
	 wire n_111;
	 wire n_109;
	 wire n_113;
	 wire n_114;
	 wire n_112;

endmodule

module omsp_alu(alu_out,alu_out_add,alu_stat,alu_stat_wr,dbg_halt_st,exec_cycle,inst_alu,inst_bw,inst_jmp,inst_so,op_dst,op_src,status);
	 output [15:0]alu_out;
	 output [15:0]alu_out_add;
	 output [3:0]alu_stat;
	 output [3:0]alu_stat_wr;
	 input dbg_halt_st;
	 input exec_cycle;
	 input [11:0]inst_alu;
	 input inst_bw;
	 input [7:0]inst_jmp;
	 input [7:0]inst_so;
	 input [15:0]op_dst;
	 input [15:0]op_src;
	 input [3:0]status;

	 wire op_bit8_msk;
	 wire op_src_inv_cmd;
	 wire n_4_0;
	 wire n_4_1;
	 wire n_4_2;
	 wire n_4_3;
	 wire n_4_4;
	 wire n_4_5;
	 wire [3:0]X;
	 wire n_4_6;
	 wire n_4_7;
	 wire n_4_8;
	 wire n_5_0;
	 wire n_5_1;
	 wire n_5_2;
	 wire n_5_3;
	 wire n_5_4;
	 wire n_5_5;
	 wire n_6_0;
	 wire alu_short_thro;
	 wire n_7_0;
	 wire n_7_1;
	 wire n_7_2;
	 wire n_7_3;
	 wire n_7_4;
	 wire n_7_5;
	 wire n_7_6;
	 wire n_7_7;
	 wire n_7_8;
	 wire n_7_9;
	 wire n_7_10;
	 wire n_7_11;
	 wire n_7_12;
	 wire n_7_13;
	 wire n_7_14;
	 wire n_7_15;
	 wire n_7_16;
	 wire n_7_17;
	 wire n_7_18;
	 wire n_7_19;
	 wire n_7_20;
	 wire n_7_21;
	 wire n_7_22;
	 wire n_7_23;
	 wire n_7_24;
	 wire n_7_25;
	 wire n_7_26;
	 wire n_7_27;
	 wire n_7_28;
	 wire n_7_29;
	 wire n_7_30;
	 wire n_7_31;
	 wire n_7_32;
	 wire n_7_33;
	 wire n_7_34;
	 wire n_7_35;
	 wire n_7_36;
	 wire n_7_37;
	 wire n_7_38;
	 wire n_7_39;
	 wire n_7_40;
	 wire n_7_41;
	 wire n_7_42;
	 wire n_7_43;
	 wire n_7_44;
	 wire n_7_45;
	 wire n_7_46;
	 wire n_7_47;
	 wire n_7_48;
	 wire n_7_49;
	 wire n_7_50;
	 wire n_7_51;
	 wire n_7_52;
	 wire n_7_53;
	 wire n_7_54;
	 wire n_7_55;
	 wire n_7_56;
	 wire n_7_57;
	 wire n_7_58;
	 wire n_7_59;
	 wire n_7_60;
	 wire n_7_61;
	 wire n_7_62;
	 wire n_7_63;
	 wire n_7_64;
	 wire n_7_65;
	 wire n_7_66;
	 wire n_7_67;
	 wire n_7_68;
	 wire n_7_69;
	 wire n_7_70;
	 wire n_7_71;
	 wire n_7_72;
	 wire n_7_73;
	 wire n_7_74;
	 wire n_7_75;
	 wire n_7_76;
	 wire n_7_77;
	 wire n_7_78;
	 wire n_7_79;
	 wire n_7_80;
	 wire n_7_81;
	 wire n_7_82;
	 wire n_7_83;
	 wire n_7_84;
	 wire n_7_85;
	 wire n_7_86;
	 wire n_7_87;
	 wire n_7_88;
	 wire n_7_89;
	 wire n_7_90;
	 wire n_7_91;
	 wire n_7_92;
	 wire n_7_93;
	 wire n_7_94;
	 wire n_7_95;
	 wire n_7_96;
	 wire n_7_97;
	 wire n_7_98;
	 wire n_7_99;
	 wire n_7_100;
	 wire n_7_101;
	 wire n_7_102;
	 wire n_7_103;
	 wire n_7_104;
	 wire n_7_105;
	 wire n_7_106;
	 wire n_7_107;
	 wire n_7_108;
	 wire n_7_109;
	 wire n_7_110;
	 wire n_7_111;
	 wire n_7_112;
	 wire n_7_113;
	 wire n_7_114;
	 wire n_7_115;
	 wire n_7_116;
	 wire n_7_117;
	 wire n_7_118;
	 wire n_7_119;
	 wire n_7_120;
	 wire n_7_121;
	 wire n_7_122;
	 wire n_7_123;
	 wire n_7_124;
	 wire n_7_125;
	 wire n_7_126;
	 wire n_7_127;
	 wire n_7_128;
	 wire n_7_129;
	 wire n_7_130;
	 wire n_7_131;
	 wire n_7_132;
	 wire n_7_133;
	 wire n_7_134;
	 wire n_7_135;
	 wire n_8_0;
	 wire n_9_0;
	 wire n_9_1;
	 wire n_9_2;
	 wire n_9_3;
	 wire n_9_4;
	 wire n_9_5;
	 wire n_9_6;
	 wire n_9_7;
	 wire n_9_8;
	 wire n_9_9;
	 wire n_11_0;
	 wire n_11_1;
	 wire n_11_2;
	 wire n_12_0;
	 wire [4:0]bcd_add;
	 wire n_12_1;
	 wire n_12_2;
	 wire n_12_3;
	 wire n_12_4;
	 wire n_12_5;
	 wire n_12_6;
	 wire n_12_7;
	 wire n_12_8;
	 wire n_13_0;
	 wire n_14_0;
	 wire n_14_1;
	 wire n_14_2;
	 wire n_14_3;
	 wire n_14_4;
	 wire n_14_5;
	 wire n_14_6;
	 wire n_14_7;
	 wire n_14_8;
	 wire n_14_9;
	 wire n_16_0;
	 wire n_16_1;
	 wire n_16_2;
	 wire n_17_0;
	 wire [4:0]bcd_add0;
	 wire n_17_1;
	 wire n_17_2;
	 wire n_17_3;
	 wire n_17_4;
	 wire n_17_5;
	 wire n_17_6;
	 wire n_17_7;
	 wire n_17_8;
	 wire n_18_0;
	 wire n_19_0;
	 wire n_19_1;
	 wire n_19_2;
	 wire n_19_3;
	 wire n_19_4;
	 wire n_19_5;
	 wire n_19_6;
	 wire n_19_7;
	 wire n_19_8;
	 wire n_19_9;
	 wire n_21_0;
	 wire n_21_1;
	 wire n_21_2;
	 wire n_22_0;
	 wire [4:0]bcd_add1;
	 wire n_22_1;
	 wire n_22_2;
	 wire n_22_3;
	 wire n_22_4;
	 wire n_22_5;
	 wire n_22_6;
	 wire n_22_7;
	 wire n_22_8;
	 wire n_23_0;
	 wire n_24_0;
	 wire n_24_1;
	 wire n_24_2;
	 wire n_24_3;
	 wire n_24_4;
	 wire n_24_5;
	 wire n_24_6;
	 wire n_24_7;
	 wire n_24_8;
	 wire n_24_9;
	 wire n_26_0;
	 wire n_26_1;
	 wire n_26_2;
	 wire n_27_0;
	 wire [4:0]bcd_add2;
	 wire n_27_1;
	 wire n_27_2;
	 wire n_27_3;
	 wire n_27_4;
	 wire n_27_5;
	 wire n_27_6;
	 wire n_27_7;
	 wire n_27_8;
	 wire n_28_0;
	 wire n_28_1;
	 wire alu_inc;
	 wire n_30_0;
	 wire n_30_1;
	 wire n_30_2;
	 wire n_30_3;
	 wire n_30_4;
	 wire n_30_5;
	 wire n_30_6;
	 wire n_30_7;
	 wire n_30_8;
	 wire n_30_9;
	 wire n_40_0;
	 wire n_40_1;
	 wire n_40_2;
	 wire n_40_3;
	 wire n_40_4;
	 wire n_40_5;
	 wire n_40_6;
	 wire n_40_7;
	 wire n_40_8;
	 wire n_40_9;
	 wire n_40_10;
	 wire n_40_11;
	 wire n_40_12;
	 wire n_40_13;
	 wire n_40_14;
	 wire [16:0]alu_add;
	 wire [16:0]alu_add_inc;
	 wire n_41_0;
	 wire n_41_1;
	 wire n_41_2;
	 wire n_41_3;
	 wire n_41_4;
	 wire n_41_5;
	 wire n_41_6;
	 wire n_41_7;
	 wire n_41_8;
	 wire n_41_9;
	 wire n_41_10;
	 wire n_41_11;
	 wire n_41_12;
	 wire n_41_13;
	 wire n_41_14;
	 wire n_41_15;
	 wire n_41_16;
	 wire n_43_0;
	 wire n_44_0;
	 wire n_44_1;
	 wire n_44_2;
	 wire n_44_3;
	 wire n_44_4;
	 wire n_44_5;
	 wire n_44_6;
	 wire n_44_7;
	 wire n_44_8;
	 wire n_44_9;
	 wire n_44_10;
	 wire n_44_11;
	 wire n_44_12;
	 wire n_44_13;
	 wire n_44_14;
	 wire n_44_15;
	 wire n_44_16;
	 wire n_46_0;
	 wire n_46_1;
	 wire n_46_2;
	 wire n_48_0;
	 wire n_48_1;
	 wire n_48_2;
	 wire n_49_0;
	 wire n_49_1;
	 wire n_49_2;
	 wire n_49_3;
	 wire n_49_4;
	 wire n_49_5;
	 wire n_49_6;
	 wire n_49_7;
	 wire n_49_8;
	 wire n_49_9;
	 wire Z;
	 wire n_51_0;
	 wire n_51_1;
	 wire n_51_2;
	 wire n_51_3;
	 wire n_51_4;
	 wire n_51_5;
	 wire n_51_6;
	 wire n_51_7;
	 wire n_51_8;
	 wire n_51_9;
	 wire n_51_10;
	 wire n_51_11;
	 wire n_51_12;
	 wire n_51_13;
	 wire n_51_14;
	 wire n_51_15;
	 wire n_51_16;
	 wire n_51_17;
	 wire n_51_18;
	 wire n_51_19;
	 wire n_51_20;
	 wire n_51_21;
	 wire n_51_22;
	 wire n_104;
	 wire n_7;
	 wire n_86;
	 wire n_87;
	 wire n_103;
	 wire n_6;
	 wire n_102;
	 wire n_5;
	 wire n_101;
	 wire n_4;
	 wire n_100;
	 wire n_3;
	 wire n_19;
	 wire n_99;
	 wire n_2;
	 wire n_18;
	 wire n_98;
	 wire n_1;
	 wire n_17;
	 wire n_97;
	 wire n_0;
	 wire n_16;
	 wire n_96;
	 wire n_15;
	 wire n_95;
	 wire n_14;
	 wire n_94;
	 wire n_13;
	 wire n_93;
	 wire n_12;
	 wire n_92;
	 wire n_11;
	 wire n_91;
	 wire n_10;
	 wire n_90;
	 wire n_9;
	 wire n_89;
	 wire n_8;
	 wire n_88;
	 wire n_106;
	 wire n_68;
	 wire n_67;
	 wire n_66;
	 wire n_65;
	 wire n_56;
	 wire n_55;
	 wire n_54;
	 wire n_53;
	 wire n_44;
	 wire n_43;
	 wire n_42;
	 wire n_41;
	 wire n_38;
	 wire n_40;
	 wire n_39;
	 wire n_45;
	 wire n_46;
	 wire n_47;
	 wire n_48;
	 wire n_49;
	 wire n_50;
	 wire n_52;
	 wire n_51;
	 wire n_57;
	 wire n_58;
	 wire n_59;
	 wire n_60;
	 wire n_61;
	 wire n_62;
	 wire n_64;
	 wire n_63;
	 wire n_69;
	 wire n_70;
	 wire n_71;
	 wire n_72;
	 wire n_73;
	 wire n_74;
	 wire n_76;
	 wire n_75;
	 wire n_78;
	 wire n_77;
	 wire n_83;
	 wire n_80;
	 wire n_79;
	 wire n_81;
	 wire n_82;
	 wire n_84;
	 wire n_105;
	 wire n_20;
	 wire n_37;
	 wire n_36;
	 wire n_35;
	 wire n_34;
	 wire n_33;
	 wire n_32;
	 wire n_31;
	 wire n_30;
	 wire n_21;
	 wire n_29;
	 wire n_28;
	 wire n_27;
	 wire n_26;
	 wire n_25;
	 wire n_24;
	 wire n_23;
	 wire n_22;
	 wire n_108;
	 wire n_110;
	 wire n_109;
	 wire n_111;
	 wire n_112;
	 wire n_85;
	 wire n_107;

	assign alu_stat_wr[3] = alu_stat_wr[0];
	assign alu_stat_wr[2] = alu_stat_wr[0];
	assign alu_stat_wr[1] = alu_stat_wr[0];
endmodule

module OAI222_X1_LVT(ZN,A1,A2,B1,B2,C1,C2);
	 output ZN;
	 input A1;
	 input A2;
	 input B1;
	 input B2;
	 input C1;
	 input C2;


endmodule

module OAI221_X1_LVT(ZN,A,B1,B2,C1,C2);
	 output ZN;
	 input A;
	 input B1;
	 input B2;
	 input C1;
	 input C2;


endmodule

module AND4_X1_LVT(ZN,A1,A2,A3,A4);
	 output ZN;
	 input A1;
	 input A2;
	 input A3;
	 input A4;


endmodule

module omsp_and_gate__2_49(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_and_gate__2_29(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_and_gate__2_47(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module openMSP430(aclk,aclk_en,dbg_freeze,dbg_i2c_sda_out,dbg_uart_txd,dco_enable,dco_wkup,dmem_addr,dmem_cen,dmem_din,dmem_wen,irq_acc,lfxt_enable,lfxt_wkup,mclk,dma_dout,dma_ready,dma_resp,per_addr,per_din,per_en,per_we,pmem_addr,pmem_cen,pmem_din,pmem_wen,puc_rst,smclk,smclk_en,cpu_en,dbg_en,dbg_i2c_addr,dbg_i2c_broadcast,dbg_i2c_scl,dbg_i2c_sda_in,dbg_uart_rxd,dco_clk,dmem_dout,irq,lfxt_clk,dma_addr,dma_din,dma_en,dma_priority,dma_we,dma_wkup,nmi,per_dout,pmem_dout,reset_n,scan_enable,scan_mode,wkup);
	 output aclk;
	 output aclk_en;
	 output dbg_freeze;
	 output dbg_i2c_sda_out;
	 output dbg_uart_txd;
	 output dco_enable;
	 output dco_wkup;
	 output [8:0]dmem_addr;
	 output dmem_cen;
	 output [15:0]dmem_din;
	 output [1:0]dmem_wen;
	 output [13:0]irq_acc;
	 output lfxt_enable;
	 output lfxt_wkup;
	 output mclk;
	 output [15:0]dma_dout;
	 output dma_ready;
	 output dma_resp;
	 output [13:0]per_addr;
	 output [15:0]per_din;
	 output per_en;
	 output [1:0]per_we;
	 output [10:0]pmem_addr;
	 output pmem_cen;
	 output [15:0]pmem_din;
	 output [1:0]pmem_wen;
	 output puc_rst;
	 output smclk;
	 output smclk_en;
	 input cpu_en;
	 input dbg_en;
	 input [6:0]dbg_i2c_addr;
	 input [6:0]dbg_i2c_broadcast;
	 input dbg_i2c_scl;
	 input dbg_i2c_sda_in;
	 input dbg_uart_rxd;
	 input dco_clk;
	 input [15:0]dmem_dout;
	 input [13:0]irq;
	 input lfxt_clk;
	 input [14:0]dma_addr;
	 input [15:0]dma_din;
	 input dma_en;
	 input dma_priority;
	 input [1:0]dma_we;
	 input dma_wkup;
	 input nmi;
	 input [15:0]per_dout;
	 input [15:0]pmem_dout;
	 input reset_n;
	 input scan_enable;
	 input scan_mode;
	 input wkup;

	 wire wdtnmies;
	 wire wdtifg;
	 wire wdt_wkup;
	 wire wdt_reset;
	 wire wdt_irq;
	 wire [15:0]per_dout_wdog;
	 wire scg1;
	 wire scg0;
	 wire pc_sw_wr;
	 wire [15:0]pc_sw;
	 wire oscoff;
	 wire [15:0]eu_mdb_out;
	 wire [1:0]eu_mb_wr;
	 wire eu_mb_en;
	 wire [15:0]eu_mab;
	 wire gie;
	 wire [15:0]dbg_reg_din;
	 wire cpuoff;
	 wire [15:0]pc_nxt;
	 wire [15:0]pc;
	 wire nmi_acc;
	 wire mclk_wkup;
	 wire mclk_enable;
	 wire mclk_dma_wkup;
	 wire mclk_dma_enable;
	 wire fe_mb_en;
	 wire [2:0]inst_type;
	 wire [15:0]inst_src;
	 wire [7:0]inst_so;
	 wire [15:0]inst_sext;
	 wire inst_mov;
	 wire [7:0]inst_jmp;
	 wire inst_irq_rst;
	 wire [15:0]inst_dext;
	 wire [15:0]inst_dest;
	 wire inst_bw;
	 wire [11:0]inst_alu;
	 wire [7:0]inst_as;
	 wire [7:0]inst_ad;
	 wire exec_done;
	 wire [3:0]e_state;
	 wire decode_noirq;
	 wire cpu_halt_st;
	 wire [15:0]per_dout_mpy;
	 wire fe_pmem_wait;
	 wire [15:0]fe_mdb_in;
	 wire [15:0]eu_mdb_in;
	 wire [15:0]dbg_mem_din;
	 wire cpu_halt_cmd;
	 wire dbg_reg_wr;
	 wire [1:0]dbg_mem_wr;
	 wire dbg_mem_en;
	 wire [15:0]dbg_mem_dout;
	 wire [15:0]dbg_mem_addr;
	 wire dbg_halt_cmd;
	 wire dbg_cpu_reset;
	 wire wdtifg_sw_set;
	 wire wdtifg_sw_clr;
	 wire wdtie;
	 wire [15:0]per_dout_sfr;
	 wire nmi_wkup;
	 wire nmi_pnd;
	 wire [31:0]cpu_id;
	 wire puc_pnd_set;
	 wire por;
	 wire [15:0]per_dout_clk;
	 wire dbg_rst;
	 wire dbg_en_s;
	 wire dbg_clk;
	 wire cpu_mclk;
	 wire cpu_en_s;
	 wire n_0_0_0;
	 wire [15:0]per_dout_or;
	 wire n_0_0_1;
	 wire n_0_0_2;
	 wire n_0_0_3;
	 wire n_0_0_4;
	 wire n_0_0_5;
	 wire n_0_0_6;
	 wire n_0_0_7;
	 wire n_0_0_8;
	 wire n_0_0_9;
	 wire n_0_0_10;
	 wire n_0_0_11;
	 wire n_0_0_12;
	 wire n_0_0_13;
	 wire n_0_0_14;
	 wire n_0_0_15;
	 wire n_14;
	 wire n_13;
	 wire n_12;
	 wire n_11;
	 wire n_10;
	 wire n_9;
	 wire n_8;
	 wire n_7;
	 wire n_6;
	 wire n_5;
	 wire n_4;
	 wire n_3;
	 wire n_2;
	 wire n_1;
	 wire n_0;
	 wire uc_0;

endmodule

module omsp_sync_cell__1_13(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_mem_backbone(cpu_halt_cmd,dbg_mem_din,dmem_addr,dmem_cen,dmem_din,dmem_wen,eu_mdb_in,fe_mdb_in,fe_pmem_wait,dma_dout,dma_ready,dma_resp,per_addr,per_din,per_we,per_en,pmem_addr,pmem_cen,pmem_din,pmem_wen,cpu_halt_st,dbg_halt_cmd,dbg_mem_addr,dbg_mem_dout,dbg_mem_en,dbg_mem_wr,dmem_dout,eu_mab,eu_mb_en,eu_mb_wr,eu_mdb_out,fe_mab,fe_mb_en,mclk,dma_addr,dma_din,dma_en,dma_priority,dma_we,per_dout,pmem_dout,puc_rst,scan_enable);
	 output cpu_halt_cmd;
	 output [15:0]dbg_mem_din;
	 output [8:0]dmem_addr;
	 output dmem_cen;
	 output [15:0]dmem_din;
	 output [1:0]dmem_wen;
	 output [15:0]eu_mdb_in;
	 output [15:0]fe_mdb_in;
	 output fe_pmem_wait;
	 output [15:0]dma_dout;
	 output dma_ready;
	 output dma_resp;
	 output [13:0]per_addr;
	 output [15:0]per_din;
	 output [1:0]per_we;
	 output per_en;
	 output [10:0]pmem_addr;
	 output pmem_cen;
	 output [15:0]pmem_din;
	 output [1:0]pmem_wen;
	 input cpu_halt_st;
	 input dbg_halt_cmd;
	 input [14:0]dbg_mem_addr;
	 input [15:0]dbg_mem_dout;
	 input dbg_mem_en;
	 input [1:0]dbg_mem_wr;
	 input [15:0]dmem_dout;
	 input [14:0]eu_mab;
	 input eu_mb_en;
	 input [1:0]eu_mb_wr;
	 input [15:0]eu_mdb_out;
	 input [14:0]fe_mab;
	 input fe_mb_en;
	 input mclk;
	 input [14:0]dma_addr;
	 input [15:0]dma_din;
	 input dma_en;
	 input dma_priority;
	 input [1:0]dma_we;
	 input [15:0]per_dout;
	 input [15:0]pmem_dout;
	 input puc_rst;
	 input scan_enable;

	 wire n_0_0;
	 wire [15:0]per_dout_val;
	 wire n_2_0;
	 wire n_2_1;
	 wire [14:0]ext_mem_addr;
	 wire n_2_2;
	 wire n_2_3;
	 wire n_2_4;
	 wire n_2_5;
	 wire n_2_6;
	 wire n_2_7;
	 wire n_2_8;
	 wire n_2_9;
	 wire n_2_10;
	 wire n_2_11;
	 wire n_2_12;
	 wire n_2_13;
	 wire n_2_14;
	 wire n_2_15;
	 wire n_3_0;
	 wire ext_per_sel;
	 wire ext_mem_en;
	 wire n_5_0;
	 wire n_5_1;
	 wire n_5_2;
	 wire eu_per_en;
	 wire n_6_0;
	 wire ext_per_en;
	 wire ext_pmem_sel;
	 wire n_8_0;
	 wire fe_pmem_en;
	 wire n_11_0;
	 wire n_11_1;
	 wire eu_pmem_en;
	 wire n_12_0;
	 wire ext_pmem_en;
	 wire [1:0]ext_mem_din_sel;
	 wire n_15_0;
	 wire n_16_0;
	 wire n_16_1;
	 wire n_16_2;
	 wire n_16_3;
	 wire n_16_4;
	 wire n_16_5;
	 wire n_16_6;
	 wire n_16_7;
	 wire n_16_8;
	 wire n_16_9;
	 wire n_16_10;
	 wire n_16_11;
	 wire n_16_12;
	 wire n_16_13;
	 wire n_16_14;
	 wire n_16_15;
	 wire n_19_0;
	 wire n_19_1;
	 wire n_19_2;
	 wire n_19_3;
	 wire n_19_4;
	 wire n_19_5;
	 wire n_19_6;
	 wire ext_dmem_sel;
	 wire n_20_0;
	 wire n_20_1;
	 wire n_20_2;
	 wire n_20_3;
	 wire n_20_4;
	 wire n_20_5;
	 wire eu_dmem_en;
	 wire n_21_0;
	 wire ext_dmem_en;
	 wire n_22_0;
	 wire n_22_1;
	 wire n_22_2;
	 wire n_22_3;
	 wire n_22_4;
	 wire n_22_5;
	 wire n_22_6;
	 wire n_22_7;
	 wire n_22_8;
	 wire n_22_9;
	 wire n_24_0;
	 wire n_24_1;
	 wire n_24_2;
	 wire n_24_3;
	 wire n_24_4;
	 wire n_24_5;
	 wire n_24_6;
	 wire n_24_7;
	 wire n_24_8;
	 wire n_24_9;
	 wire n_24_10;
	 wire n_24_11;
	 wire n_24_12;
	 wire n_24_13;
	 wire n_24_14;
	 wire n_24_15;
	 wire n_24_16;
	 wire n_25_0;
	 wire n_25_1;
	 wire n_25_2;
	 wire n_25_3;
	 wire n_25_4;
	 wire n_25_5;
	 wire n_25_6;
	 wire n_25_7;
	 wire n_25_8;
	 wire n_25_9;
	 wire n_25_10;
	 wire n_25_11;
	 wire n_25_12;
	 wire n_25_13;
	 wire n_25_14;
	 wire n_25_15;
	 wire n_25_16;
	 wire n_27_0;
	 wire n_27_1;
	 wire [1:0]ext_mem_wr;
	 wire n_27_2;
	 wire n_29_0;
	 wire n_29_1;
	 wire n_29_2;
	 wire [1:0]eu_mdb_in_sel;
	 wire n_31_0;
	 wire n_32_0;
	 wire n_32_1;
	 wire n_32_2;
	 wire n_32_3;
	 wire n_32_4;
	 wire n_32_5;
	 wire n_32_6;
	 wire n_32_7;
	 wire n_32_8;
	 wire n_32_9;
	 wire n_32_10;
	 wire n_32_11;
	 wire n_32_12;
	 wire n_32_13;
	 wire n_32_14;
	 wire n_32_15;
	 wire fe_pmem_en_dly;
	 wire n_33_0;
	 wire fe_pmem_save;
	 wire [15:0]pmem_dout_bckup;
	 wire n_35_0;
	 wire n_35_1;
	 wire fe_pmem_restore;
	 wire pmem_dout_bckup_sel;
	 wire n_37_0;
	 wire n_37_1;
	 wire n_39_0;
	 wire n_39_1;
	 wire n_39_2;
	 wire n_39_3;
	 wire n_39_4;
	 wire n_39_5;
	 wire n_39_6;
	 wire n_39_7;
	 wire n_39_8;
	 wire n_39_9;
	 wire n_39_10;
	 wire n_39_11;
	 wire n_39_12;
	 wire n_39_13;
	 wire n_39_14;
	 wire n_39_15;
	 wire n_39_16;
	 wire n_42_0;
	 wire n_43_0;
	 wire dma_ready_dly;
	 wire n_45_0;
	 wire n_45_1;
	 wire n_45_2;
	 wire n_45_3;
	 wire n_45_4;
	 wire n_45_5;
	 wire n_45_6;
	 wire n_45_7;
	 wire n_45_8;
	 wire n_46_0;
	 wire n_46_1;
	 wire n_46_2;
	 wire n_46_3;
	 wire n_46_4;
	 wire n_46_5;
	 wire n_46_6;
	 wire n_46_7;
	 wire n_46_8;
	 wire n_46_9;
	 wire n_46_10;
	 wire n_46_11;
	 wire n_46_12;
	 wire n_46_13;
	 wire n_46_14;
	 wire n_46_15;
	 wire n_46_16;
	 wire n_47_0;
	 wire n_47_1;
	 wire n_47_2;
	 wire n_49_0;
	 wire n_49_1;
	 wire n_49_2;
	 wire n_49_3;
	 wire n_49_4;
	 wire n_49_5;
	 wire n_49_6;
	 wire n_49_7;
	 wire n_49_8;
	 wire n_49_9;
	 wire n_49_10;
	 wire n_49_11;
	 wire n_51_0;
	 wire n_51_1;
	 wire n_0;
	 wire n_1;
	 wire n_2;
	 wire n_4;
	 wire n_3;
	 wire n_5;
	 wire n_6;
	 wire n_8;
	 wire n_10;
	 wire n_7;
	 wire n_9;
	 wire n_12;
	 wire n_11;
	 wire n_15;
	 wire n_14;
	 wire n_13;
	 wire n_16;

	assign per_addr[8] = 1'b0;
	assign per_addr[9] = 1'b1;
	assign per_addr[10] = 1'b2;
	assign per_addr[11] = 1'b3;
	assign per_addr[12] = 1'b4;
	assign per_addr[13] = 1'b5;
endmodule

module omsp_register_file(cpuoff,gie,oscoff,pc_sw,pc_sw_wr,reg_dest,reg_src,scg0,scg1,status,alu_stat,alu_stat_wr,inst_bw,inst_dest,inst_src,mclk,pc,puc_rst,reg_dest_val,reg_dest_wr,reg_pc_call,reg_sp_val,reg_sp_wr,reg_sr_wr,reg_sr_clr,reg_incr,scan_enable);
	 output cpuoff;
	 output gie;
	 output oscoff;
	 output [15:0]pc_sw;
	 output pc_sw_wr;
	 output [15:0]reg_dest;
	 output [15:0]reg_src;
	 output scg0;
	 output scg1;
	 output [3:0]status;
	 input [3:0]alu_stat;
	 input [3:0]alu_stat_wr;
	 input inst_bw;
	 input [15:0]inst_dest;
	 input [15:0]inst_src;
	 input mclk;
	 input [15:0]pc;
	 input puc_rst;
	 input [15:0]reg_dest_val;
	 input reg_dest_wr;
	 input reg_pc_call;
	 input [15:0]reg_sp_val;
	 input reg_sp_wr;
	 input reg_sr_wr;
	 input reg_sr_clr;
	 input reg_incr;
	 input scan_enable;

	 wire n_0_0;
	 wire n_1_0;
	 wire r2_wr;
	 wire n_2_0;
	 wire n_2_1;
	 wire [4:0]r2_nxt;
	 wire n_2_2;
	 wire n_2_3;
	 wire n_2_4;
	 wire n_5_0;
	 wire n_5_1;
	 wire n_5_2;
	 wire n_5_3;
	 wire n_5_4;
	 wire n_5_5;
	 wire n_5_6;
	 wire n_5_7;
	 wire n_5_8;
	 wire n_5_9;
	 wire n_5_10;
	 wire n_5_11;
	 wire n_5_12;
	 wire n_5_13;
	 wire n_5_14;
	 wire n_5_15;
	 wire n_5_16;
	 wire n_6_0;
	 wire n_8_0;
	 wire n_9_0;
	 wire n_10_0;
	 wire inst_src_in;
	 wire r1_inc;
	 wire r1_wr;
	 wire n_13_0;
	 wire n_13_1;
	 wire n_14_0;
	 wire r3_wr;
	 wire [15:0]r3;
	 wire n_17_0;
	 wire r4_inc;
	 wire r4_wr;
	 wire n_20_0;
	 wire [15:0]reg_incr_val;
	 wire n_22_0;
	 wire n_22_1;
	 wire n_22_2;
	 wire n_22_3;
	 wire n_22_4;
	 wire n_22_5;
	 wire n_22_6;
	 wire n_22_7;
	 wire n_22_8;
	 wire n_22_9;
	 wire n_22_10;
	 wire n_22_11;
	 wire n_22_12;
	 wire n_22_13;
	 wire n_22_14;
	 wire n_22_15;
	 wire [15:0]r4;
	 wire n_24_0;
	 wire n_24_1;
	 wire n_24_2;
	 wire n_24_3;
	 wire n_24_4;
	 wire n_24_5;
	 wire n_24_6;
	 wire n_24_7;
	 wire n_24_8;
	 wire n_24_9;
	 wire n_24_10;
	 wire n_24_11;
	 wire n_24_12;
	 wire n_24_13;
	 wire n_24_14;
	 wire n_24_15;
	 wire n_24_16;
	 wire n_25_0;
	 wire n_25_1;
	 wire n_27_0;
	 wire r5_inc;
	 wire r5_wr;
	 wire [15:0]r5;
	 wire n_31_0;
	 wire n_31_1;
	 wire n_31_2;
	 wire n_31_3;
	 wire n_31_4;
	 wire n_31_5;
	 wire n_31_6;
	 wire n_31_7;
	 wire n_31_8;
	 wire n_31_9;
	 wire n_31_10;
	 wire n_31_11;
	 wire n_31_12;
	 wire n_31_13;
	 wire n_31_14;
	 wire n_31_15;
	 wire n_31_16;
	 wire n_32_0;
	 wire n_32_1;
	 wire n_34_0;
	 wire r6_inc;
	 wire r6_wr;
	 wire [15:0]r6;
	 wire n_38_0;
	 wire n_38_1;
	 wire n_38_2;
	 wire n_38_3;
	 wire n_38_4;
	 wire n_38_5;
	 wire n_38_6;
	 wire n_38_7;
	 wire n_38_8;
	 wire n_38_9;
	 wire n_38_10;
	 wire n_38_11;
	 wire n_38_12;
	 wire n_38_13;
	 wire n_38_14;
	 wire n_38_15;
	 wire n_38_16;
	 wire n_39_0;
	 wire n_39_1;
	 wire n_41_0;
	 wire r7_inc;
	 wire r7_wr;
	 wire [15:0]r7;
	 wire n_45_0;
	 wire n_45_1;
	 wire n_45_2;
	 wire n_45_3;
	 wire n_45_4;
	 wire n_45_5;
	 wire n_45_6;
	 wire n_45_7;
	 wire n_45_8;
	 wire n_45_9;
	 wire n_45_10;
	 wire n_45_11;
	 wire n_45_12;
	 wire n_45_13;
	 wire n_45_14;
	 wire n_45_15;
	 wire n_45_16;
	 wire n_46_0;
	 wire n_46_1;
	 wire n_48_0;
	 wire r8_inc;
	 wire r8_wr;
	 wire [15:0]r8;
	 wire n_52_0;
	 wire n_52_1;
	 wire n_52_2;
	 wire n_52_3;
	 wire n_52_4;
	 wire n_52_5;
	 wire n_52_6;
	 wire n_52_7;
	 wire n_52_8;
	 wire n_52_9;
	 wire n_52_10;
	 wire n_52_11;
	 wire n_52_12;
	 wire n_52_13;
	 wire n_52_14;
	 wire n_52_15;
	 wire n_52_16;
	 wire n_53_0;
	 wire n_53_1;
	 wire n_55_0;
	 wire r9_inc;
	 wire r9_wr;
	 wire [15:0]r9;
	 wire n_59_0;
	 wire n_59_1;
	 wire n_59_2;
	 wire n_59_3;
	 wire n_59_4;
	 wire n_59_5;
	 wire n_59_6;
	 wire n_59_7;
	 wire n_59_8;
	 wire n_59_9;
	 wire n_59_10;
	 wire n_59_11;
	 wire n_59_12;
	 wire n_59_13;
	 wire n_59_14;
	 wire n_59_15;
	 wire n_59_16;
	 wire n_60_0;
	 wire n_60_1;
	 wire n_62_0;
	 wire r10_inc;
	 wire r10_wr;
	 wire [15:0]r10;
	 wire n_66_0;
	 wire n_66_1;
	 wire n_66_2;
	 wire n_66_3;
	 wire n_66_4;
	 wire n_66_5;
	 wire n_66_6;
	 wire n_66_7;
	 wire n_66_8;
	 wire n_66_9;
	 wire n_66_10;
	 wire n_66_11;
	 wire n_66_12;
	 wire n_66_13;
	 wire n_66_14;
	 wire n_66_15;
	 wire n_66_16;
	 wire n_67_0;
	 wire n_67_1;
	 wire n_69_0;
	 wire r11_inc;
	 wire r11_wr;
	 wire [15:0]r11;
	 wire n_73_0;
	 wire n_73_1;
	 wire n_73_2;
	 wire n_73_3;
	 wire n_73_4;
	 wire n_73_5;
	 wire n_73_6;
	 wire n_73_7;
	 wire n_73_8;
	 wire n_73_9;
	 wire n_73_10;
	 wire n_73_11;
	 wire n_73_12;
	 wire n_73_13;
	 wire n_73_14;
	 wire n_73_15;
	 wire n_73_16;
	 wire n_74_0;
	 wire n_74_1;
	 wire n_76_0;
	 wire r12_inc;
	 wire r12_wr;
	 wire [15:0]r12;
	 wire n_80_0;
	 wire n_80_1;
	 wire n_80_2;
	 wire n_80_3;
	 wire n_80_4;
	 wire n_80_5;
	 wire n_80_6;
	 wire n_80_7;
	 wire n_80_8;
	 wire n_80_9;
	 wire n_80_10;
	 wire n_80_11;
	 wire n_80_12;
	 wire n_80_13;
	 wire n_80_14;
	 wire n_80_15;
	 wire n_80_16;
	 wire n_81_0;
	 wire n_81_1;
	 wire n_83_0;
	 wire r13_inc;
	 wire r13_wr;
	 wire [15:0]r13;
	 wire n_87_0;
	 wire n_87_1;
	 wire n_87_2;
	 wire n_87_3;
	 wire n_87_4;
	 wire n_87_5;
	 wire n_87_6;
	 wire n_87_7;
	 wire n_87_8;
	 wire n_87_9;
	 wire n_87_10;
	 wire n_87_11;
	 wire n_87_12;
	 wire n_87_13;
	 wire n_87_14;
	 wire n_87_15;
	 wire n_87_16;
	 wire n_88_0;
	 wire n_88_1;
	 wire n_90_0;
	 wire r14_inc;
	 wire r14_wr;
	 wire [15:0]r14;
	 wire n_94_0;
	 wire n_94_1;
	 wire n_94_2;
	 wire n_94_3;
	 wire n_94_4;
	 wire n_94_5;
	 wire n_94_6;
	 wire n_94_7;
	 wire n_94_8;
	 wire n_94_9;
	 wire n_94_10;
	 wire n_94_11;
	 wire n_94_12;
	 wire n_94_13;
	 wire n_94_14;
	 wire n_94_15;
	 wire n_94_16;
	 wire n_95_0;
	 wire n_95_1;
	 wire n_97_0;
	 wire r15_inc;
	 wire r15_wr;
	 wire [15:0]r15;
	 wire n_101_0;
	 wire n_101_1;
	 wire n_101_2;
	 wire n_101_3;
	 wire n_101_4;
	 wire n_101_5;
	 wire n_101_6;
	 wire n_101_7;
	 wire n_101_8;
	 wire n_101_9;
	 wire n_101_10;
	 wire n_101_11;
	 wire n_101_12;
	 wire n_101_13;
	 wire n_101_14;
	 wire n_101_15;
	 wire n_101_16;
	 wire n_102_0;
	 wire n_102_1;
	 wire n_104_0;
	 wire n_105_0;
	 wire n_105_1;
	 wire n_105_2;
	 wire n_105_3;
	 wire n_105_4;
	 wire n_105_5;
	 wire n_105_6;
	 wire n_105_7;
	 wire n_105_8;
	 wire n_105_9;
	 wire n_105_10;
	 wire n_105_11;
	 wire n_105_12;
	 wire n_105_13;
	 wire n_105_14;
	 wire n_105_15;
	 wire n_105_16;
	 wire n_105_17;
	 wire n_105_18;
	 wire n_105_19;
	 wire n_105_20;
	 wire n_105_21;
	 wire n_105_22;
	 wire n_105_23;
	 wire n_105_24;
	 wire n_105_25;
	 wire n_105_26;
	 wire n_105_27;
	 wire n_105_28;
	 wire n_105_29;
	 wire n_105_30;
	 wire n_105_31;
	 wire n_105_32;
	 wire n_105_33;
	 wire n_105_34;
	 wire n_105_35;
	 wire n_105_36;
	 wire n_105_37;
	 wire n_105_38;
	 wire n_105_39;
	 wire n_105_40;
	 wire n_105_41;
	 wire n_105_42;
	 wire n_105_43;
	 wire n_105_44;
	 wire n_105_45;
	 wire n_105_46;
	 wire n_105_47;
	 wire n_105_48;
	 wire n_105_49;
	 wire n_105_50;
	 wire n_105_51;
	 wire n_105_52;
	 wire n_105_53;
	 wire n_105_54;
	 wire n_105_55;
	 wire n_105_56;
	 wire n_105_57;
	 wire n_105_58;
	 wire n_105_59;
	 wire n_105_60;
	 wire n_105_61;
	 wire n_105_62;
	 wire n_105_63;
	 wire n_105_64;
	 wire n_105_65;
	 wire n_105_66;
	 wire n_105_67;
	 wire n_105_68;
	 wire n_105_69;
	 wire n_105_70;
	 wire n_105_71;
	 wire n_105_72;
	 wire n_105_73;
	 wire n_105_74;
	 wire n_105_75;
	 wire n_105_76;
	 wire n_105_77;
	 wire n_105_78;
	 wire n_105_79;
	 wire n_105_80;
	 wire n_105_81;
	 wire n_105_82;
	 wire n_105_83;
	 wire n_105_84;
	 wire n_105_85;
	 wire n_105_86;
	 wire n_105_87;
	 wire n_105_88;
	 wire n_105_89;
	 wire n_105_90;
	 wire n_105_91;
	 wire n_105_92;
	 wire n_105_93;
	 wire n_105_94;
	 wire n_105_95;
	 wire n_105_96;
	 wire n_105_97;
	 wire n_105_98;
	 wire n_105_99;
	 wire n_105_100;
	 wire n_105_101;
	 wire n_105_102;
	 wire n_105_103;
	 wire n_105_104;
	 wire n_105_105;
	 wire n_105_106;
	 wire n_105_107;
	 wire n_105_108;
	 wire n_105_109;
	 wire n_105_110;
	 wire n_105_111;
	 wire n_105_112;
	 wire n_105_113;
	 wire n_105_114;
	 wire n_105_115;
	 wire n_105_116;
	 wire n_105_117;
	 wire n_105_118;
	 wire n_105_119;
	 wire n_105_120;
	 wire n_105_121;
	 wire n_105_122;
	 wire n_105_123;
	 wire n_105_124;
	 wire n_105_125;
	 wire n_105_126;
	 wire n_105_127;
	 wire n_105_128;
	 wire n_105_129;
	 wire n_105_130;
	 wire n_105_131;
	 wire n_105_132;
	 wire n_105_133;
	 wire n_105_134;
	 wire n_105_135;
	 wire n_105_136;
	 wire n_105_137;
	 wire n_105_138;
	 wire n_105_139;
	 wire n_105_140;
	 wire n_105_141;
	 wire n_105_142;
	 wire n_105_143;
	 wire n_105_144;
	 wire n_105_145;
	 wire n_105_146;
	 wire n_105_147;
	 wire n_105_148;
	 wire n_105_149;
	 wire n_105_150;
	 wire n_105_151;
	 wire n_105_152;
	 wire n_105_153;
	 wire n_105_154;
	 wire n_105_155;
	 wire n_105_156;
	 wire n_105_157;
	 wire n_105_158;
	 wire n_105_159;
	 wire n_105_160;
	 wire n_105_161;
	 wire n_105_162;
	 wire n_105_163;
	 wire n_105_164;
	 wire n_105_165;
	 wire n_105_166;
	 wire n_105_167;
	 wire n_105_168;
	 wire n_105_169;
	 wire n_105_170;
	 wire n_105_171;
	 wire n_105_172;
	 wire n_105_173;
	 wire n_105_174;
	 wire n_105_175;
	 wire n_105_176;
	 wire n_105_177;
	 wire n_105_178;
	 wire n_105_179;
	 wire n_105_180;
	 wire n_105_181;
	 wire n_105_182;
	 wire n_105_183;
	 wire n_105_184;
	 wire n_105_185;
	 wire n_105_186;
	 wire n_105_187;
	 wire n_105_188;
	 wire n_105_189;
	 wire n_105_190;
	 wire n_105_191;
	 wire n_105_192;
	 wire n_105_193;
	 wire n_105_194;
	 wire n_105_195;
	 wire n_105_196;
	 wire n_105_197;
	 wire n_105_198;
	 wire n_105_199;
	 wire n_105_200;
	 wire n_105_201;
	 wire n_105_202;
	 wire n_105_203;
	 wire n_105_204;
	 wire n_105_205;
	 wire n_105_206;
	 wire n_105_207;
	 wire n_105_208;
	 wire n_105_209;
	 wire n_105_210;
	 wire n_105_211;
	 wire n_105_212;
	 wire n_105_213;
	 wire n_105_214;
	 wire n_105_215;
	 wire n_105_216;
	 wire n_105_217;
	 wire n_105_218;
	 wire n_105_219;
	 wire n_105_220;
	 wire n_105_221;
	 wire n_105_222;
	 wire n_105_223;
	 wire n_105_224;
	 wire n_105_225;
	 wire n_105_226;
	 wire n_105_227;
	 wire n_105_228;
	 wire n_105_229;
	 wire n_105_230;
	 wire n_105_231;
	 wire n_105_232;
	 wire n_105_233;
	 wire n_105_234;
	 wire n_105_235;
	 wire n_105_236;
	 wire n_105_237;
	 wire n_105_238;
	 wire n_105_239;
	 wire n_105_240;
	 wire n_105_241;
	 wire n_105_242;
	 wire n_105_243;
	 wire n_105_244;
	 wire n_105_245;
	 wire n_105_246;
	 wire n_105_247;
	 wire n_105_248;
	 wire n_105_249;
	 wire n_105_250;
	 wire n_105_251;
	 wire n_105_252;
	 wire n_105_253;
	 wire n_105_254;
	 wire n_105_255;
	 wire n_105_256;
	 wire n_105_257;
	 wire n_105_258;
	 wire n_105_259;
	 wire n_105_260;
	 wire n_105_261;
	 wire n_105_262;
	 wire n_105_263;
	 wire n_105_264;
	 wire n_105_265;
	 wire n_105_266;
	 wire n_105_267;
	 wire n_105_268;
	 wire n_105_269;
	 wire n_105_270;
	 wire n_105_271;
	 wire n_105_272;
	 wire n_105_273;
	 wire n_105_274;
	 wire n_105_275;
	 wire n_105_276;
	 wire n_105_277;
	 wire n_105_278;
	 wire n_105_279;
	 wire n_105_280;
	 wire n_105_281;
	 wire n_105_282;
	 wire n_105_283;
	 wire n_105_284;
	 wire n_105_285;
	 wire n_105_286;
	 wire n_105_287;
	 wire n_105_288;
	 wire n_105_289;
	 wire n_105_290;
	 wire n_105_291;
	 wire n_105_292;
	 wire n_105_293;
	 wire n_105_294;
	 wire n_105_295;
	 wire n_105_296;
	 wire n_105_297;
	 wire n_105_298;
	 wire n_105_299;
	 wire n_105_300;
	 wire n_105_301;
	 wire n_105_302;
	 wire n_105_303;
	 wire n_105_304;
	 wire n_105_305;
	 wire n_105_306;
	 wire n_105_307;
	 wire n_105_308;
	 wire n_105_309;
	 wire n_105_310;
	 wire n_105_311;
	 wire n_105_312;
	 wire n_105_313;
	 wire n_105_314;
	 wire n_105_315;
	 wire n_105_316;
	 wire n_105_317;
	 wire n_105_318;
	 wire n_105_319;
	 wire n_106_0;
	 wire n_106_1;
	 wire n_106_2;
	 wire n_106_3;
	 wire n_106_4;
	 wire n_106_5;
	 wire n_106_6;
	 wire n_106_7;
	 wire n_106_8;
	 wire n_106_9;
	 wire n_106_10;
	 wire n_106_11;
	 wire n_106_12;
	 wire n_106_13;
	 wire [15:0]r1;
	 wire n_108_0;
	 wire n_109_0;
	 wire n_109_1;
	 wire n_109_2;
	 wire n_109_3;
	 wire n_109_4;
	 wire n_109_5;
	 wire n_109_6;
	 wire n_109_7;
	 wire n_109_8;
	 wire n_109_9;
	 wire n_109_10;
	 wire n_109_11;
	 wire n_109_12;
	 wire n_109_13;
	 wire n_109_14;
	 wire n_110_0;
	 wire n_110_1;
	 wire n_110_2;
	 wire n_112_0;
	 wire n_112_1;
	 wire n_112_2;
	 wire n_112_3;
	 wire n_112_4;
	 wire n_112_5;
	 wire n_112_6;
	 wire n_112_7;
	 wire n_112_8;
	 wire n_112_9;
	 wire n_112_10;
	 wire n_112_11;
	 wire n_112_12;
	 wire n_112_13;
	 wire n_112_14;
	 wire n_112_15;
	 wire n_112_16;
	 wire n_112_17;
	 wire n_112_18;
	 wire n_112_19;
	 wire n_112_20;
	 wire n_112_21;
	 wire n_112_22;
	 wire n_112_23;
	 wire n_112_24;
	 wire n_112_25;
	 wire n_112_26;
	 wire n_112_27;
	 wire n_112_28;
	 wire n_112_29;
	 wire n_112_30;
	 wire n_112_31;
	 wire n_112_32;
	 wire n_112_33;
	 wire n_112_34;
	 wire n_112_35;
	 wire n_112_36;
	 wire n_112_37;
	 wire n_112_38;
	 wire n_112_39;
	 wire n_112_40;
	 wire n_112_41;
	 wire n_112_42;
	 wire n_112_43;
	 wire n_112_44;
	 wire n_112_45;
	 wire n_112_46;
	 wire n_112_47;
	 wire n_112_48;
	 wire n_112_49;
	 wire n_112_50;
	 wire n_112_51;
	 wire n_112_52;
	 wire n_112_53;
	 wire n_112_54;
	 wire n_112_55;
	 wire n_112_56;
	 wire n_112_57;
	 wire n_112_58;
	 wire n_112_59;
	 wire n_112_60;
	 wire n_112_61;
	 wire n_112_62;
	 wire n_112_63;
	 wire n_112_64;
	 wire n_112_65;
	 wire n_112_66;
	 wire n_112_67;
	 wire n_112_68;
	 wire n_112_69;
	 wire n_112_70;
	 wire n_112_71;
	 wire n_112_72;
	 wire n_112_73;
	 wire n_112_74;
	 wire n_112_75;
	 wire n_112_76;
	 wire n_112_77;
	 wire n_112_78;
	 wire n_112_79;
	 wire n_112_80;
	 wire n_112_81;
	 wire n_112_82;
	 wire n_112_83;
	 wire n_112_84;
	 wire n_112_85;
	 wire n_112_86;
	 wire n_112_87;
	 wire n_112_88;
	 wire n_112_89;
	 wire n_112_90;
	 wire n_112_91;
	 wire n_112_92;
	 wire n_112_93;
	 wire n_112_94;
	 wire n_112_95;
	 wire n_112_96;
	 wire n_112_97;
	 wire n_112_98;
	 wire n_112_99;
	 wire n_112_100;
	 wire n_112_101;
	 wire n_112_102;
	 wire n_112_103;
	 wire n_112_104;
	 wire n_112_105;
	 wire n_112_106;
	 wire n_112_107;
	 wire n_112_108;
	 wire n_112_109;
	 wire n_112_110;
	 wire n_112_111;
	 wire n_112_112;
	 wire n_112_113;
	 wire n_112_114;
	 wire n_112_115;
	 wire n_112_116;
	 wire n_112_117;
	 wire n_112_118;
	 wire n_112_119;
	 wire n_112_120;
	 wire n_112_121;
	 wire n_112_122;
	 wire n_112_123;
	 wire n_112_124;
	 wire n_112_125;
	 wire n_112_126;
	 wire n_112_127;
	 wire n_112_128;
	 wire n_112_129;
	 wire n_112_130;
	 wire n_112_131;
	 wire n_112_132;
	 wire n_112_133;
	 wire n_112_134;
	 wire n_112_135;
	 wire n_112_136;
	 wire n_112_137;
	 wire n_112_138;
	 wire n_112_139;
	 wire n_112_140;
	 wire n_112_141;
	 wire n_112_142;
	 wire n_112_143;
	 wire n_112_144;
	 wire n_112_145;
	 wire n_112_146;
	 wire n_112_147;
	 wire n_112_148;
	 wire n_112_149;
	 wire n_112_150;
	 wire n_112_151;
	 wire n_112_152;
	 wire n_112_153;
	 wire n_112_154;
	 wire n_112_155;
	 wire n_112_156;
	 wire n_112_157;
	 wire n_112_158;
	 wire n_112_159;
	 wire n_112_160;
	 wire n_112_161;
	 wire n_112_162;
	 wire n_112_163;
	 wire n_112_164;
	 wire n_112_165;
	 wire n_112_166;
	 wire n_112_167;
	 wire n_112_168;
	 wire n_112_169;
	 wire n_112_170;
	 wire n_112_171;
	 wire n_112_172;
	 wire n_112_173;
	 wire n_112_174;
	 wire n_112_175;
	 wire n_112_176;
	 wire n_112_177;
	 wire n_112_178;
	 wire n_112_179;
	 wire n_112_180;
	 wire n_112_181;
	 wire n_112_182;
	 wire n_112_183;
	 wire n_112_184;
	 wire n_112_185;
	 wire n_112_186;
	 wire n_112_187;
	 wire n_112_188;
	 wire n_112_189;
	 wire n_112_190;
	 wire n_112_191;
	 wire n_112_192;
	 wire n_112_193;
	 wire n_112_194;
	 wire n_112_195;
	 wire n_112_196;
	 wire n_112_197;
	 wire n_112_198;
	 wire n_112_199;
	 wire n_112_200;
	 wire n_112_201;
	 wire n_112_202;
	 wire n_112_203;
	 wire n_112_204;
	 wire n_112_205;
	 wire n_112_206;
	 wire n_112_207;
	 wire n_112_208;
	 wire n_112_209;
	 wire n_112_210;
	 wire n_112_211;
	 wire n_112_212;
	 wire n_112_213;
	 wire n_112_214;
	 wire n_112_215;
	 wire n_112_216;
	 wire n_112_217;
	 wire n_112_218;
	 wire n_112_219;
	 wire n_112_220;
	 wire n_112_221;
	 wire n_112_222;
	 wire n_112_223;
	 wire n_112_224;
	 wire n_112_225;
	 wire n_112_226;
	 wire n_112_227;
	 wire n_112_228;
	 wire n_112_229;
	 wire n_112_230;
	 wire n_112_231;
	 wire n_112_232;
	 wire n_112_233;
	 wire n_112_234;
	 wire n_112_235;
	 wire n_112_236;
	 wire n_112_237;
	 wire n_112_238;
	 wire n_112_239;
	 wire n_112_240;
	 wire n_112_241;
	 wire n_112_242;
	 wire n_112_243;
	 wire n_112_244;
	 wire n_112_245;
	 wire n_112_246;
	 wire n_112_247;
	 wire n_112_248;
	 wire n_112_249;
	 wire n_112_250;
	 wire n_112_251;
	 wire n_112_252;
	 wire n_112_253;
	 wire n_112_254;
	 wire n_112_255;
	 wire n_112_256;
	 wire n_112_257;
	 wire n_112_258;
	 wire n_112_259;
	 wire n_112_260;
	 wire n_112_261;
	 wire n_112_262;
	 wire n_112_263;
	 wire n_112_264;
	 wire n_112_265;
	 wire n_112_266;
	 wire n_112_267;
	 wire n_112_268;
	 wire n_112_269;
	 wire n_112_270;
	 wire n_112_271;
	 wire n_112_272;
	 wire n_112_273;
	 wire n_112_274;
	 wire n_112_275;
	 wire n_112_276;
	 wire n_112_277;
	 wire n_112_278;
	 wire n_112_279;
	 wire n_112_280;
	 wire n_112_281;
	 wire n_112_282;
	 wire n_112_283;
	 wire n_112_284;
	 wire n_112_285;
	 wire n_112_286;
	 wire n_112_287;
	 wire n_112_288;
	 wire n_112_289;
	 wire n_112_290;
	 wire n_112_291;
	 wire n_112_292;
	 wire n_112_293;
	 wire n_112_294;
	 wire n_112_295;
	 wire n_112_296;
	 wire n_112_297;
	 wire n_112_298;
	 wire n_112_299;
	 wire n_112_300;
	 wire n_112_301;
	 wire n_112_302;
	 wire n_112_303;
	 wire n_112_304;
	 wire n_112_305;
	 wire n_112_306;
	 wire n_112_307;
	 wire n_112_308;
	 wire n_112_309;
	 wire n_112_310;
	 wire n_112_311;
	 wire n_112_312;
	 wire n_112_313;
	 wire n_112_314;
	 wire n_112_315;
	 wire n_112_316;
	 wire n_112_317;
	 wire n_112_318;
	 wire n_112_319;
	 wire n_7;
	 wire n_17;
	 wire n_8;
	 wire n_16;
	 wire n_24;
	 wire n_22;
	 wire n_23;
	 wire n_21;
	 wire n_0;
	 wire n_272;
	 wire n_271;
	 wire n_41;
	 wire n_44;
	 wire n_27;
	 wire n_2;
	 wire n_39;
	 wire n_4;
	 wire n_37;
	 wire n_6;
	 wire n_35;
	 wire n_19;
	 wire n_33;
	 wire n_31;
	 wire n_25;
	 wire n_26;
	 wire n_29;
	 wire n_10;
	 wire n_14;
	 wire n_255;
	 wire n_273;
	 wire n_288;
	 wire n_270;
	 wire n_178;
	 wire n_181;
	 wire n_196;
	 wire n_179;
	 wire n_159;
	 wire n_162;
	 wire n_177;
	 wire n_160;
	 wire n_140;
	 wire n_143;
	 wire n_158;
	 wire n_141;
	 wire n_121;
	 wire n_124;
	 wire n_139;
	 wire n_122;
	 wire n_102;
	 wire n_105;
	 wire n_120;
	 wire n_103;
	 wire n_83;
	 wire n_86;
	 wire n_101;
	 wire n_84;
	 wire n_64;
	 wire n_67;
	 wire n_82;
	 wire n_65;
	 wire n_45;
	 wire n_48;
	 wire n_63;
	 wire n_46;
	 wire n_197;
	 wire n_200;
	 wire n_215;
	 wire n_198;
	 wire n_254;
	 wire n_235;
	 wire n_238;
	 wire n_253;
	 wire n_236;
	 wire n_216;
	 wire n_219;
	 wire n_234;
	 wire n_217;
	 wire n_28;
	 wire n_9;
	 wire n_13;
	 wire n_180;
	 wire n_161;
	 wire n_142;
	 wire n_123;
	 wire n_104;
	 wire n_85;
	 wire n_66;
	 wire n_47;
	 wire n_199;
	 wire n_237;
	 wire n_218;
	 wire n_30;
	 wire n_11;
	 wire n_15;
	 wire n_256;
	 wire n_274;
	 wire n_182;
	 wire n_163;
	 wire n_144;
	 wire n_125;
	 wire n_106;
	 wire n_87;
	 wire n_68;
	 wire n_49;
	 wire n_201;
	 wire n_239;
	 wire n_220;
	 wire n_257;
	 wire n_275;
	 wire n_183;
	 wire n_164;
	 wire n_145;
	 wire n_126;
	 wire n_107;
	 wire n_88;
	 wire n_69;
	 wire n_50;
	 wire n_202;
	 wire n_240;
	 wire n_221;
	 wire n_32;
	 wire n_258;
	 wire n_276;
	 wire n_184;
	 wire n_165;
	 wire n_146;
	 wire n_127;
	 wire n_108;
	 wire n_89;
	 wire n_70;
	 wire n_51;
	 wire n_203;
	 wire n_241;
	 wire n_222;
	 wire n_259;
	 wire n_277;
	 wire n_185;
	 wire n_166;
	 wire n_147;
	 wire n_128;
	 wire n_109;
	 wire n_90;
	 wire n_71;
	 wire n_52;
	 wire n_204;
	 wire n_242;
	 wire n_223;
	 wire n_34;
	 wire n_18;
	 wire n_260;
	 wire n_278;
	 wire n_186;
	 wire n_167;
	 wire n_148;
	 wire n_129;
	 wire n_110;
	 wire n_91;
	 wire n_72;
	 wire n_53;
	 wire n_205;
	 wire n_243;
	 wire n_224;
	 wire n_261;
	 wire n_279;
	 wire n_187;
	 wire n_168;
	 wire n_149;
	 wire n_130;
	 wire n_111;
	 wire n_92;
	 wire n_73;
	 wire n_54;
	 wire n_206;
	 wire n_244;
	 wire n_225;
	 wire n_36;
	 wire n_12;
	 wire n_20;
	 wire n_262;
	 wire n_280;
	 wire n_188;
	 wire n_169;
	 wire n_150;
	 wire n_131;
	 wire n_112;
	 wire n_93;
	 wire n_74;
	 wire n_55;
	 wire n_207;
	 wire n_245;
	 wire n_226;
	 wire n_263;
	 wire n_281;
	 wire n_189;
	 wire n_170;
	 wire n_151;
	 wire n_132;
	 wire n_113;
	 wire n_94;
	 wire n_75;
	 wire n_56;
	 wire n_208;
	 wire n_246;
	 wire n_227;
	 wire n_38;
	 wire n_5;
	 wire n_264;
	 wire n_282;
	 wire n_190;
	 wire n_171;
	 wire n_152;
	 wire n_133;
	 wire n_114;
	 wire n_95;
	 wire n_76;
	 wire n_57;
	 wire n_209;
	 wire n_247;
	 wire n_228;
	 wire n_265;
	 wire n_283;
	 wire n_191;
	 wire n_172;
	 wire n_153;
	 wire n_134;
	 wire n_115;
	 wire n_96;
	 wire n_77;
	 wire n_58;
	 wire n_210;
	 wire n_248;
	 wire n_229;
	 wire n_40;
	 wire n_3;
	 wire n_266;
	 wire n_284;
	 wire n_192;
	 wire n_173;
	 wire n_154;
	 wire n_135;
	 wire n_116;
	 wire n_97;
	 wire n_78;
	 wire n_59;
	 wire n_211;
	 wire n_249;
	 wire n_230;
	 wire n_267;
	 wire n_285;
	 wire n_193;
	 wire n_174;
	 wire n_155;
	 wire n_136;
	 wire n_117;
	 wire n_98;
	 wire n_79;
	 wire n_60;
	 wire n_212;
	 wire n_250;
	 wire n_231;
	 wire n_42;
	 wire n_1;
	 wire n_268;
	 wire n_286;
	 wire n_194;
	 wire n_175;
	 wire n_156;
	 wire n_137;
	 wire n_118;
	 wire n_99;
	 wire n_80;
	 wire n_61;
	 wire n_213;
	 wire n_251;
	 wire n_232;
	 wire n_269;
	 wire n_287;
	 wire n_195;
	 wire n_176;
	 wire n_157;
	 wire n_138;
	 wire n_119;
	 wire n_100;
	 wire n_81;
	 wire n_62;
	 wire n_214;
	 wire n_252;
	 wire n_233;
	 wire n_43;

	assign pc_sw[0] = reg_dest_val[0];
	assign pc_sw[1] = reg_dest_val[1];
	assign pc_sw[2] = reg_dest_val[2];
	assign pc_sw[3] = reg_dest_val[3];
	assign pc_sw[4] = reg_dest_val[4];
	assign pc_sw[5] = reg_dest_val[5];
	assign pc_sw[6] = reg_dest_val[6];
	assign pc_sw[7] = reg_dest_val[7];
endmodule

module omsp_and_gate__2_35(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_sync_cell__2_19(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_clock_gate__2_3(gclk,clk,enable,scan_enable);
	 output gclk;
	 input clk;
	 input enable;
	 input scan_enable;

	 wire enable_in;
	 wire enable_latch;
	 wire n_0;

endmodule

module omsp_scan_mux__1_9(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module omsp_clock_gate__2_7(gclk,clk,enable,scan_enable);
	 output gclk;
	 input clk;
	 input enable;
	 input scan_enable;

	 wire enable_in;
	 wire enable_latch;
	 wire n_0;

endmodule

module OR3_X1_LVT(ZN,A1,A2,A3);
	 output ZN;
	 input A1;
	 input A2;
	 input A3;


endmodule

module omsp_sync_reset__0_1432(rst_s,clk,rst_a);
	 output rst_s;
	 input clk;
	 input rst_a;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_clock_gate__2_15(gclk,clk,enable,scan_enable);
	 output gclk;
	 input clk;
	 input enable;
	 input scan_enable;

	 wire enable_in;
	 wire enable_latch;
	 wire n_0;

endmodule

module omsp_sync_reset(rst_s,clk,rst_a);
	 output rst_s;
	 input clk;
	 input rst_a;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_and_gate__2_37(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_scan_mux__2_61(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module omsp_and_gate__2_31(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_clock_gate__2_11(gclk,clk,enable,scan_enable);
	 output gclk;
	 input clk;
	 input enable;
	 input scan_enable;

	 wire enable_in;
	 wire enable_latch;
	 wire n_0;

endmodule

module XOR2_X1_LVT(Z,A,B);
	 output Z;
	 input A;
	 input B;


endmodule

module NOR2_X1_LVT(ZN,A1,A2);
	 output ZN;
	 input A1;
	 input A2;


endmodule

module omsp_scan_mux__1_7(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module omsp_scan_mux__2_65(data_out,data_in_scan,data_in_func,scan_mode);
	 output data_out;
	 input data_in_scan;
	 input data_in_func;
	 input scan_mode;

	 wire n_0_0;
	 wire n_0_1;

endmodule

module omsp_and_gate__2_45(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_sync_cell__2_25(data_out,clk,data_in,rst);
	 output data_out;
	 input clk;
	 input data_in;
	 input rst;

	 wire n_0;
	 wire n_1;

endmodule

module omsp_and_gate__2_51(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_wakeup_cell(wkup_out,scan_clk,scan_mode,scan_rst,wkup_clear,wkup_event);
	 output wkup_out;
	 input scan_clk;
	 input scan_mode;
	 input scan_rst;
	 input wkup_clear;
	 input wkup_event;

	 wire wkup_rst;
	 wire wkup_clk;
	 wire n_0;

endmodule

module omsp_and_gate__2_33(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

module omsp_and_gate__2_39(y,a,b);
	 output y;
	 input a;
	 input b;


endmodule

