`celldefine

module ADDFXL (S, CO, A, B, CI);
output S, CO;
input A, B, CI;
endmodule

module ADDFX1 (S, CO, A, B, CI);
output S, CO;
input A, B, CI;
endmodule

module ADDFX2 (S, CO, A, B, CI);
output S, CO;
input A, B, CI;
endmodule

module ADDFX4 (S, CO, A, B, CI);
output S, CO;
input A, B, CI;
endmodule

module ADDFHXL (S, CO, A, B, CI);
output S, CO;
input A, B, CI;
endmodule

module ADDFHX1 (S, CO, A, B, CI);
output S, CO;
input A, B, CI;
endmodule

module ADDFHX2 (S, CO, A, B, CI);
output S, CO;
input A, B, CI;
endmodule

module ADDFHX4 (S, CO, A, B, CI);
output S, CO;
input A, B, CI;
endmodule

module ADDHXL (S, CO, A, B);
output S, CO;
input A, B;
endmodule

module ADDHX1 (S, CO, A, B);
output S, CO;
input A, B;
endmodule

module ADDHX2 (S, CO, A, B);
output S, CO;
input A, B;
endmodule

module ADDHX4 (S, CO, A, B);
output S, CO;
input A, B;
endmodule

module AND2XL (Y, A, B);
output Y;
input A, B;
endmodule

module AND2X1 (Y, A, B);
output Y;
input A, B;
endmodule

module AND2X2 (Y, A, B);
output Y;
input A, B;
endmodule

module AND2X4 (Y, A, B);
output Y;
input A, B;
endmodule

module AND3XL (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module AND3X1 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module AND3X2 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module AND3X4 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module AND4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module AND4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module AND4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module AND4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module AOI21XL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;
endmodule

module AOI21X1 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;
endmodule

module AOI21X2 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;
endmodule

module AOI21X4 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;
endmodule

module AOI211XL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;
endmodule

module AOI211X1 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;
endmodule

module AOI211X2 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;
endmodule

module AOI211X4 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;
endmodule

module AOI22XL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;
endmodule

module AOI22X1 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;
endmodule

module AOI22X2 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;
endmodule

module AOI22X4 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;
endmodule

module AOI221XL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;
endmodule

module AOI221X1 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;
endmodule

module AOI221X2 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;
endmodule

module AOI221X4 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;
endmodule

module AOI222XL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;
endmodule

module AOI222X1 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;
endmodule

module AOI222X2 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;
endmodule

module AOI222X4 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;
endmodule

module AOI2BB1XL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;
endmodule

module AOI2BB1X1 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;
endmodule

module AOI2BB1X2 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;
endmodule

module AOI2BB1X4 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;
endmodule

module AOI2BB2XL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;
endmodule

module AOI2BB2X1 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;
endmodule

module AOI2BB2X2 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;
endmodule

module AOI2BB2X4 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;
endmodule

module AOI31XL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;
endmodule

module AOI31X1 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;
endmodule

module AOI31X2 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;
endmodule

module AOI31X4 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;
endmodule

module AOI32XL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;
endmodule

module AOI32X1 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;
endmodule

module AOI32X2 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;
endmodule

module AOI32X4 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;
endmodule

module AOI33XL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;
endmodule

module AOI33X1 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;
endmodule

module AOI33X2 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;
endmodule

module AOI33X4 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;
endmodule

module BUFXL (Y, A);
output Y;
input A;
endmodule

module BUFX1 (Y, A);
output Y;
input A;
endmodule

module BUFX2 (Y, A);
output Y;
input A;
endmodule

module BUFX3 (Y, A);
output Y;
input A;
endmodule

module BUFX4 (Y, A);
output Y;
input A;
endmodule

module BUFX8 (Y, A);
output Y;
input A;
endmodule

module BUFX12 (Y, A);
output Y;
input A;
endmodule

module BUFX16 (Y, A);
output Y;
input A;
endmodule

module BUFX20 (Y, A);
output Y;
input A;
endmodule

module CLKBUFXL (Y, A);
output Y;
input A;
endmodule

module CLKBUFX1 (Y, A);
output Y;
input A;
endmodule

module CLKBUFX2 (Y, A);
output Y;
input A;
endmodule

module CLKBUFX3 (Y, A);
output Y;
input A;
endmodule

module CLKBUFX4 (Y, A);
output Y;
input A;
endmodule

module CLKBUFX8 (Y, A);
output Y;
input A;
endmodule

module CLKBUFX12 (Y, A);
output Y;
input A;
endmodule

module CLKBUFX16 (Y, A);
output Y;
input A;
endmodule

module CLKBUFX20 (Y, A);
output Y;
input A;
endmodule

module CLKINVXL (Y, A);
output Y;
input A;
endmodule

module CLKINVX1 (Y, A);
output Y;
input A;
endmodule

module CLKINVX2 (Y, A);
output Y;
input A;
endmodule

module CLKINVX3 (Y, A);
output Y;
input A;
endmodule

module CLKINVX4 (Y, A);
output Y;
input A;
endmodule

module CLKINVX8 (Y, A);
output Y;
input A;
endmodule

module CLKINVX12 (Y, A);
output Y;
input A;
endmodule

module CLKINVX16 (Y, A);
output Y;
input A;
endmodule

module CLKINVX20 (Y, A);
output Y;
input A;
endmodule

module JKFFXL (Q, QN, J, K, CK);
output Q, QN;
input J, K, CK;
endmodule

module JKFFX1 (Q, QN, J, K, CK);
output Q, QN;
input J, K, CK;
endmodule

module JKFFX2 (Q, QN, J, K, CK);
output Q, QN;
input J, K, CK;
endmodule

module JKFFX4 (Q, QN, J, K, CK);
output Q, QN;
input J, K, CK;
endmodule

module JKFFRXL (Q, QN, J, K, CK, RN);
output Q, QN;
input J, K, CK, RN;
endmodule

module JKFFRX1 (Q, QN, J, K, CK, RN);
output Q, QN;
input J, K, CK, RN;
endmodule

module JKFFRX2 (Q, QN, J, K, CK, RN);
output Q, QN;
input J, K, CK, RN;
endmodule

module JKFFRX4 (Q, QN, J, K, CK, RN);
output Q, QN;
input J, K, CK, RN;
endmodule

module JKFFSXL (Q, QN, J, K, CK, SN);
output Q, QN;
input J, K, CK, SN;
endmodule

module JKFFSX1 (Q, QN, J, K, CK, SN);
output Q, QN;
input J, K, CK, SN;
endmodule

module JKFFSX2 (Q, QN, J, K, CK, SN);
output Q, QN;
input J, K, CK, SN;
endmodule

module JKFFSX4 (Q, QN, J, K, CK, SN);
output Q, QN;
input J, K, CK, SN;
endmodule

module JKFFSRXL (Q, QN, J, K, CK, SN, RN);
output Q, QN;
input J, K, CK, SN, RN;
endmodule

module JKFFSRX1 (Q, QN, J, K, CK, SN, RN);
output Q, QN;
input J, K, CK, SN, RN;
endmodule

module JKFFSRX2 (Q, QN, J, K, CK, SN, RN);
output Q, QN;
input J, K, CK, SN, RN;
endmodule

module JKFFSRX4 (Q, QN, J, K, CK, SN, RN);
output Q, QN;
input J, K, CK, SN, RN;
endmodule

module DFFXL (Q, QN, D, CK);
output Q, QN;
input D, CK;
endmodule

module DFFX1 (Q, QN, D, CK);
output Q, QN;
input D, CK;
endmodule

module DFFX2 (Q, QN, D, CK);
output Q, QN;
input D, CK;
endmodule

module DFFX4 (Q, QN, D, CK);
output Q, QN;
input D, CK;
endmodule

module DFFHQXL (Q, D, CK);
output Q;
input D, CK;
endmodule

module DFFHQX1 (Q, D, CK);
output Q;
input D, CK;
endmodule

module DFFHQX2 (Q, D, CK);
output Q;
input D, CK;
endmodule

module DFFHQX4 (Q, D, CK);
output Q;
input D, CK;
endmodule

module DFFNSRXL (Q, QN, D, CKN, SN, RN);
output Q, QN;
input D, CKN, SN, RN;
endmodule

module DFFNSRX1 (Q, QN, D, CKN, SN, RN);
output Q, QN;
input D, CKN, SN, RN;
endmodule

module DFFNSRX2 (Q, QN, D, CKN, SN, RN);
output Q, QN;
input D, CKN, SN, RN;
endmodule

module DFFNSRX4 (Q, QN, D, CKN, SN, RN);
output Q, QN;
input D, CKN, SN, RN;
endmodule

module DFFRXL (Q, QN, D, CK, RN);
output Q, QN;
input D, CK, RN;
endmodule

module DFFRX1 (Q, QN, D, CK, RN);
output Q, QN;
input D, CK, RN;
endmodule

module DFFRX2 (Q, QN, D, CK, RN);
output Q, QN;
input D, CK, RN;
endmodule

module DFFRX4 (Q, QN, D, CK, RN);
output Q, QN;
input D, CK, RN;
endmodule

module DFFRHQXL (Q, D, CK, RN);
output Q;
input D, CK, RN;
endmodule

module DFFRHQX1 (Q, D, CK, RN);
output Q;
input D, CK, RN;
endmodule

module DFFRHQX2 (Q, D, CK, RN);
output Q;
input D, CK, RN;
endmodule

module DFFRHQX4 (Q, D, CK, RN);
output Q;
input D, CK, RN;
endmodule

module DFFSXL (Q, QN, D, CK, SN);
output Q, QN;
input D, CK, SN;
endmodule

module DFFSX1 (Q, QN, D, CK, SN);
output Q, QN;
input D, CK, SN;
endmodule

module DFFSX2 (Q, QN, D, CK, SN);
output Q, QN;
input D, CK, SN;
endmodule

module DFFSX4 (Q, QN, D, CK, SN);
output Q, QN;
input D, CK, SN;
endmodule

module DFFSHQXL (Q, D, CK, SN);
output Q;
input D, CK, SN;
endmodule

module DFFSHQX1 (Q, D, CK, SN);
output Q;
input D, CK, SN;
endmodule

module DFFSHQX2 (Q, D, CK, SN);
output Q;
input D, CK, SN;
endmodule

module DFFSHQX4 (Q, D, CK, SN);
output Q;
input D, CK, SN;
endmodule

module DFFSRXL (Q, QN, D, CK, SN, RN);
output Q, QN;
input D, CK, SN, RN;
endmodule

module DFFSRX1 (Q, QN, D, CK, SN, RN);
output Q, QN;
input D, CK, SN, RN;
endmodule

module DFFSRX2 (Q, QN, D, CK, SN, RN);
output Q, QN;
input D, CK, SN, RN;
endmodule

module DFFSRX4 (Q, QN, D, CK, SN, RN);
output Q, QN;
input D, CK, SN, RN;
endmodule

module DFFSRHQXL (Q, D, CK, SN, RN);
output Q;
input D, CK, SN, RN;
endmodule

module DFFSRHQX1 (Q, D, CK, SN, RN);
output Q;
input D, CK, SN, RN;
endmodule

module DFFSRHQX2 (Q, D, CK, SN, RN);
output Q;
input D, CK, SN, RN;
endmodule

module DFFSRHQX4 (Q, D, CK, SN, RN);
output Q;
input D, CK, SN, RN;
endmodule

module DFFTRXL (Q, QN, D, CK, RN);
output Q, QN;
input D, CK, RN;
endmodule

module DFFTRX1 (Q, QN, D, CK, RN);
output Q, QN;
input D, CK, RN;
endmodule

module DFFTRX2 (Q, QN, D, CK, RN);
output Q, QN;
input D, CK, RN;
endmodule

module DFFTRX4 (Q, QN, D, CK, RN);
output Q, QN;
input D, CK, RN;
endmodule

module DLY1X1 (Y, A);
output Y;
input A;
endmodule

module DLY2X1 (Y, A);
output Y;
input A;
endmodule

module DLY3X1 (Y, A);
output Y;
input A;
endmodule

module DLY4X1 (Y, A);
output Y;
input A;
endmodule

module EDFFXL (Q, QN, D, CK, E);
output Q, QN;
input D, CK, E;
endmodule

module EDFFX1 (Q, QN, D, CK, E);
output Q, QN;
input D, CK, E;
endmodule

module EDFFX2 (Q, QN, D, CK, E);
output Q, QN;
input D, CK, E;
endmodule

module EDFFX4 (Q, QN, D, CK, E);
output Q, QN;
input D, CK, E;
endmodule

module EDFFTRXL (Q, QN, D, CK, E, RN);
output Q, QN;
input D, CK, E, RN;
endmodule

module EDFFTRX1 (Q, QN, D, CK, E, RN);
output Q, QN;
input D, CK, E, RN;
endmodule

module EDFFTRX2 (Q, QN, D, CK, E, RN);
output Q, QN;
input D, CK, E, RN;
endmodule

module EDFFTRX4 (Q, QN, D, CK, E, RN);
output Q, QN;
input D, CK, E, RN;
endmodule

module INVXL (Y, A);
output Y;
input A;
endmodule

module INVX1 (Y, A);
output Y;
input A;
endmodule

module INVX2 (Y, A);
output Y;
input A;
endmodule

module INVX3 (Y, A);
output Y;
input A;
endmodule

module INVX4 (Y, A);
output Y;
input A;
endmodule

module INVX8 (Y, A);
output Y;
input A;
endmodule

module INVX12 (Y, A);
output Y;
input A;
endmodule

module INVX16 (Y, A);
output Y;
input A;
endmodule

module INVX20 (Y, A);
output Y;
input A;
endmodule

module MX2XL (Y, A, B, S0);
output Y;
input A, B, S0;
endmodule

module MX2X1 (Y, A, B, S0);
output Y;
input A, B, S0;
endmodule

module MX2X2 (Y, A, B, S0);
output Y;
input A, B, S0;
endmodule

module MX2X4 (Y, A, B, S0);
output Y;
input A, B, S0;
endmodule

module MX4XL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;
endmodule

module MX4X1 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;
endmodule

module MX4X2 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;
endmodule

module MX4X4 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;
endmodule

module MXI2XL (Y, A, B, S0);
output Y;
input A, B, S0;
endmodule

module MXI2X1 (Y, A, B, S0);
output Y;
input A, B, S0;
endmodule

module MXI2X2 (Y, A, B, S0);
output Y;
input A, B, S0;
endmodule

module MXI2X4 (Y, A, B, S0);
output Y;
input A, B, S0;
endmodule

module MXI4XL (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;
endmodule

module MXI4X1 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;
endmodule

module MXI4X2 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;
endmodule

module MXI4X4 (Y, A, B, C, D, S0, S1);
output Y;
input A, B, C, D, S0, S1;
endmodule

module NAND2XL (Y, A, B);
output Y;
input A, B;
endmodule

module NAND2X1 (Y, A, B);
output Y;
input A, B;
endmodule

module NAND2X2 (Y, A, B);
output Y;
input A, B;
endmodule

module NAND2X4 (Y, A, B);
output Y;
input A, B;
endmodule

module NAND2BXL (Y, AN, B);
output Y;
input AN, B;
endmodule

module NAND2BX1 (Y, AN, B);
output Y;
input AN, B;
endmodule

module NAND2BX2 (Y, AN, B);
output Y;
input AN, B;
endmodule

module NAND2BX4 (Y, AN, B);
output Y;
input AN, B;
endmodule

module NAND3XL (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module NAND3X1 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module NAND3X2 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module NAND3X4 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module NAND3BXL (Y, AN, B, C);
output Y;
input AN, B, C;
endmodule

module NAND3BX1 (Y, AN, B, C);
output Y;
input AN, B, C;
endmodule

module NAND3BX2 (Y, AN, B, C);
output Y;
input AN, B, C;
endmodule

module NAND3BX4 (Y, AN, B, C);
output Y;
input AN, B, C;
endmodule

module NAND4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module NAND4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module NAND4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module NAND4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module NAND4BXL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;
endmodule

module NAND4BX1 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;
endmodule

module NAND4BX2 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;
endmodule

module NAND4BX4 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;
endmodule

module NAND4BBXL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;
endmodule

module NAND4BBX1 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;
endmodule

module NAND4BBX2 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;
endmodule

module NAND4BBX4 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;
endmodule

module NOR2XL (Y, A, B);
output Y;
input A, B;
endmodule

module NOR2X1 (Y, A, B);
output Y;
input A, B;
endmodule

module NOR2X2 (Y, A, B);
output Y;
input A, B;
endmodule

module NOR2X4 (Y, A, B);
output Y;
input A, B;
endmodule

module NOR2BXL (Y, AN, B);
output Y;
input AN, B;
endmodule

module NOR2BX1 (Y, AN, B);
output Y;
input AN, B;
endmodule

module NOR2BX2 (Y, AN, B);
output Y;
input AN, B;
endmodule

module NOR2BX4 (Y, AN, B);
output Y;
input AN, B;
endmodule

module NOR3XL (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module NOR3X1 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module NOR3X2 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module NOR3X4 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module NOR3BXL (Y, AN, B, C);
output Y;
input AN, B, C;
endmodule

module NOR3BX1 (Y, AN, B, C);
output Y;
input AN, B, C;
endmodule

module NOR3BX2 (Y, AN, B, C);
output Y;
input AN, B, C;
endmodule

module NOR3BX4 (Y, AN, B, C);
output Y;
input AN, B, C;
endmodule

module NOR4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module NOR4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module NOR4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module NOR4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module NOR4BXL (Y, AN, B, C, D);
output Y;
input AN, B, C, D;
endmodule

module NOR4BX1 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;
endmodule

module NOR4BX2 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;
endmodule

module NOR4BX4 (Y, AN, B, C, D);
output Y;
input AN, B, C, D;
endmodule

module NOR4BBXL (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;
endmodule

module NOR4BBX1 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;
endmodule

module NOR4BBX2 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;
endmodule

module NOR4BBX4 (Y, AN, BN, C, D);
output Y;
input AN, BN, C, D;
endmodule

module OAI21XL (Y, A0, A1, B0);
output Y;
input A0, A1, B0;
endmodule

module OAI21X1 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;
endmodule

module OAI21X2 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;
endmodule

module OAI21X4 (Y, A0, A1, B0);
output Y;
input A0, A1, B0;
endmodule

module OAI211XL (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;
endmodule

module OAI211X1 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;
endmodule

module OAI211X2 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;
endmodule

module OAI211X4 (Y, A0, A1, B0, C0);
output Y;
input A0, A1, B0, C0;
endmodule

module OAI22XL (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;
endmodule

module OAI22X1 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;
endmodule

module OAI22X2 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;
endmodule

module OAI22X4 (Y, A0, A1, B0, B1);
output Y;
input A0, A1, B0, B1;
endmodule

module OAI221XL (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;
endmodule

module OAI221X1 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;
endmodule

module OAI221X2 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;
endmodule

module OAI221X4 (Y, A0, A1, B0, B1, C0);
output Y;
input A0, A1, B0, B1, C0;
endmodule

module OAI222XL (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;
endmodule

module OAI222X1 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;
endmodule

module OAI222X2 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;
endmodule

module OAI222X4 (Y, A0, A1, B0, B1, C0, C1);
output Y;
input A0, A1, B0, B1, C0, C1;
endmodule

module OAI2BB1XL (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;
endmodule

module OAI2BB1X1 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;
endmodule

module OAI2BB1X2 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;
endmodule

module OAI2BB1X4 (Y, A0N, A1N, B0);
output Y;
input A0N, A1N, B0;
endmodule

module OAI2BB2XL (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;
endmodule

module OAI2BB2X1 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;
endmodule

module OAI2BB2X2 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;
endmodule

module OAI2BB2X4 (Y, A0N, A1N, B0, B1);
output Y;
input A0N, A1N, B0, B1;
endmodule

module OAI31XL (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;
endmodule

module OAI31X1 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;
endmodule

module OAI31X2 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;
endmodule

module OAI31X4 (Y, A0, A1, A2, B0);
output Y;
input A0, A1, A2, B0;
endmodule

module OAI32XL (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;
endmodule

module OAI32X1 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;
endmodule

module OAI32X2 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;
endmodule

module OAI32X4 (Y, A0, A1, A2, B0, B1);
output Y;
input A0, A1, A2, B0, B1;
endmodule

module OAI33XL (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;
endmodule

module OAI33X1 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;
endmodule

module OAI33X2 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;
endmodule

module OAI33X4 (Y, A0, A1, A2, B0, B1, B2);
output Y;
input A0, A1, A2, B0, B1, B2;
endmodule

module OR2XL (Y, A, B);
output Y;
input A, B;
endmodule

module OR2X1 (Y, A, B);
output Y;
input A, B;
endmodule

module OR2X2 (Y, A, B);
output Y;
input A, B;
endmodule

module OR2X4 (Y, A, B);
output Y;
input A, B;
endmodule

module OR3XL (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module OR3X1 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module OR3X2 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module OR3X4 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module OR4XL (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module OR4X1 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module OR4X2 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module OR4X4 (Y, A, B, C, D);
output Y;
input A, B, C, D;
endmodule

module RSLATNXL (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
endmodule

module RSLATNX1 (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
endmodule

module RSLATNX2 (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
endmodule

module RSLATNX4 (Q, QN, RN, SN);
output Q, QN;
input RN, SN;
endmodule

module SDFFXL (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
endmodule

module SDFFX1 (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
endmodule

module SDFFX2 (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
endmodule

module SDFFX4 (Q, QN, D, SI, SE, CK);
output Q, QN;
input D, SI, SE, CK;
endmodule

module SDFFHQXL (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
endmodule

module SDFFHQX1 (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
endmodule

module SDFFHQX2 (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
endmodule

module SDFFHQX4 (Q, D, SI, SE, CK);
output Q;
input D, SI, SE, CK;
endmodule

module SDFFNSRXL (Q, QN, D, SI, SE, CKN, SN, RN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
endmodule

module SDFFNSRX1 (Q, QN, D, SI, SE, CKN, SN, RN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
endmodule

module SDFFNSRX2 (Q, QN, D, SI, SE, CKN, SN, RN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
endmodule

module SDFFNSRX4 (Q, QN, D, SI, SE, CKN, SN, RN);
output Q, QN;
input D, SI, SE, CKN, SN, RN;
endmodule

module SDFFRXL (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
endmodule

module SDFFRX1 (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
endmodule

module SDFFRX2 (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
endmodule

module SDFFRX4 (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
endmodule

module SDFFRHQXL (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
endmodule

module SDFFRHQX1 (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
endmodule

module SDFFRHQX2 (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
endmodule

module SDFFRHQX4 (Q, D, SI, SE, CK, RN);
output Q;
input D, SI, SE, CK, RN;
endmodule

module SDFFSXL (Q, QN, D, SI, SE, CK, SN);
output Q, QN;
input D, SI, SE, CK, SN;
endmodule

module SDFFSX1 (Q, QN, D, SI, SE, CK, SN);
output Q, QN;
input D, SI, SE, CK, SN;
endmodule

module SDFFSX2 (Q, QN, D, SI, SE, CK, SN);
output Q, QN;
input D, SI, SE, CK, SN;
endmodule

module SDFFSX4 (Q, QN, D, SI, SE, CK, SN);
output Q, QN;
input D, SI, SE, CK, SN;
endmodule

module SDFFSHQXL (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
endmodule

module SDFFSHQX1 (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
endmodule

module SDFFSHQX2 (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
endmodule

module SDFFSHQX4 (Q, D, SI, SE, CK, SN);
output Q;
input D, SI, SE, CK, SN;
endmodule

module SDFFSRXL (Q, QN, D, SI, SE, CK, SN, RN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
endmodule

module SDFFSRX1 (Q, QN, D, SI, SE, CK, SN, RN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
endmodule

module SDFFSRX2 (Q, QN, D, SI, SE, CK, SN, RN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
endmodule

module SDFFSRX4 (Q, QN, D, SI, SE, CK, SN, RN);
output Q, QN;
input D, SI, SE, CK, SN, RN;
endmodule

module SDFFSRHQXL (Q, D, SI, SE, CK, SN, RN);
output Q;
input D, SI, SE, CK, SN, RN;
endmodule

module SDFFSRHQX1 (Q, D, SI, SE, CK, SN, RN);
output Q;
input D, SI, SE, CK, SN, RN;
endmodule

module SDFFSRHQX2 (Q, D, SI, SE, CK, SN, RN);
output Q;
input D, SI, SE, CK, SN, RN;
endmodule

module SDFFSRHQX4 (Q, D, SI, SE, CK, SN, RN);
output Q;
input D, SI, SE, CK, SN, RN;
endmodule

module SDFFTRXL (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
endmodule

module SDFFTRX1 (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
endmodule

module SDFFTRX2 (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
endmodule

module SDFFTRX4 (Q, QN, D, SI, SE, CK, RN);
output Q, QN;
input D, SI, SE, CK, RN;
endmodule

module SEDFFXL (Q, QN, D, CK, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
endmodule

module SEDFFX1 (Q, QN, D, CK, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
endmodule

module SEDFFX2 (Q, QN, D, CK, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
endmodule

module SEDFFX4 (Q, QN, D, CK, E, SE, SI);
output Q, QN;
input D, CK, E, SE, SI;
endmodule

module SEDFFHQXL (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
endmodule

module SEDFFHQX1 (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
endmodule

module SEDFFHQX2 (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
endmodule

module SEDFFHQX4 (Q, D, CK, E, SE, SI);
output Q;
input D, CK, E, SE, SI;
endmodule

module SEDFFTRXL (Q, QN, D, CK, E, SE, SI, RN);
output Q, QN;
input D, CK, E, SE, SI, RN;
endmodule

module SEDFFTRX1 (Q, QN, D, CK, E, SE, SI, RN);
output Q, QN;
input D, CK, E, SE, SI, RN;
endmodule

module SEDFFTRX2 (Q, QN, D, CK, E, SE, SI, RN);
output Q, QN;
input D, CK, E, SE, SI, RN;
endmodule

module SEDFFTRX4 (Q, QN, D, CK, E, SE, SI, RN);
output Q, QN;
input D, CK, E, SE, SI, RN;
endmodule

module TBUFXL (Y, A, OE);
output Y;
input A, OE;
endmodule

module TBUFX1 (Y, A, OE);
output Y;
input A, OE;
endmodule

module TBUFX2 (Y, A, OE);
output Y;
input A, OE;
endmodule

module TBUFX3 (Y, A, OE);
output Y;
input A, OE;
endmodule

module TBUFX4 (Y, A, OE);
output Y;
input A, OE;
endmodule

module TBUFX8 (Y, A, OE);
output Y;
input A, OE;
endmodule

module TBUFX12 (Y, A, OE);
output Y;
input A, OE;
endmodule

module TBUFX16 (Y, A, OE);
output Y;
input A, OE;
endmodule

module TBUFX20 (Y, A, OE);
output Y;
input A, OE;
endmodule

module TIEHI (Y);
output Y;
endmodule

module TIELO (Y);
output Y;
endmodule

module TLATXL (Q, QN, D, G);
output Q, QN;
input D, G;
endmodule

module TLATX1 (Q, QN, D, G);
output Q, QN;
input D, G;
endmodule

module TLATX2 (Q, QN, D, G);
output Q, QN;
input D, G;
endmodule

module TLATX4 (Q, QN, D, G);
output Q, QN;
input D, G;
endmodule

module TLATNXL (Q, QN, D, GN);
output Q, QN;
input D, GN;
endmodule

module TLATNX1 (Q, QN, D, GN);
output Q, QN;
input D, GN;
endmodule

module TLATNX2 (Q, QN, D, GN);
output Q, QN;
input D, GN;
endmodule

module TLATNX4 (Q, QN, D, GN);
output Q, QN;
input D, GN;
endmodule

module TLATNSRXL (Q, QN, D, GN, RN, SN);
output Q, QN;
input D, GN, RN, SN;
endmodule

module TLATNSRX1 (Q, QN, D, GN, RN, SN);
output Q, QN;
input D, GN, RN, SN;
endmodule

module TLATNSRX2 (Q, QN, D, GN, RN, SN);
output Q, QN;
input D, GN, RN, SN;
endmodule

module TLATNSRX4 (Q, QN, D, GN, RN, SN);
output Q, QN;
input D, GN, RN, SN;
endmodule

module TLATSRXL (Q, QN, D, G, RN, SN);
output Q, QN;
input D, G, RN, SN;
endmodule

module TLATSRX1 (Q, QN, D, G, RN, SN);
output Q, QN;
input D, G, RN, SN;
endmodule

module TLATSRX2 (Q, QN, D, G, RN, SN);
output Q, QN;
input D, G, RN, SN;
endmodule

module TLATSRX4 (Q, QN, D, G, RN, SN);
output Q, QN;
input D, G, RN, SN;
endmodule

module XNOR2XL (Y, A, B);
output Y;
input A, B;
endmodule

module XNOR2X1 (Y, A, B);
output Y;
input A, B;
endmodule

module XNOR2X2 (Y, A, B);
output Y;
input A, B;
endmodule

module XNOR2X4 (Y, A, B);
output Y;
input A, B;
endmodule

module XNOR3X2 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module XNOR3X4 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module XOR2XL (Y, A, B);
output Y;
input A, B;
endmodule

module XOR2X1 (Y, A, B);
output Y;
input A, B;
endmodule

module XOR2X2 (Y, A, B);
output Y;
input A, B;
endmodule

module XOR2X4 (Y, A, B);
output Y;
input A, B;
endmodule

module XOR3X2 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

module XOR3X4 (Y, A, B, C);
output Y;
input A, B, C;
endmodule

`endcelldefine
